magic
tech sky130A
magscale 1 2
timestamp 1667805946
<< metal1 >>
rect 102042 700748 102048 700800
rect 102100 700788 102106 700800
rect 105446 700788 105452 700800
rect 102100 700760 105452 700788
rect 102100 700748 102106 700760
rect 105446 700748 105452 700760
rect 105504 700748 105510 700800
rect 200022 700748 200028 700800
rect 200080 700788 200086 700800
rect 202782 700788 202788 700800
rect 200080 700760 202788 700788
rect 200080 700748 200086 700760
rect 202782 700748 202788 700760
rect 202840 700748 202846 700800
rect 314470 700748 314476 700800
rect 314528 700788 314534 700800
rect 316310 700788 316316 700800
rect 314528 700760 316316 700788
rect 314528 700748 314534 700760
rect 316310 700748 316316 700760
rect 316368 700748 316374 700800
rect 53006 700544 53012 700596
rect 53064 700584 53070 700596
rect 56778 700584 56784 700596
rect 53064 700556 56784 700584
rect 53064 700544 53070 700556
rect 56778 700544 56784 700556
rect 56836 700544 56842 700596
rect 151078 700544 151084 700596
rect 151136 700584 151142 700596
rect 154114 700584 154120 700596
rect 151136 700556 154120 700584
rect 151136 700544 151142 700556
rect 154114 700544 154120 700556
rect 154172 700544 154178 700596
rect 412450 700408 412456 700460
rect 412508 700448 412514 700460
rect 413646 700448 413652 700460
rect 412508 700420 413652 700448
rect 412508 700408 412514 700420
rect 413646 700408 413652 700420
rect 413704 700408 413710 700460
rect 363506 700340 363512 700392
rect 363564 700380 363570 700392
rect 364978 700380 364984 700392
rect 363564 700352 364984 700380
rect 363564 700340 363570 700352
rect 364978 700340 364984 700352
rect 365036 700340 365042 700392
rect 20346 700204 20352 700256
rect 20404 700244 20410 700256
rect 24302 700244 24308 700256
rect 20404 700216 24308 700244
rect 20404 700204 20410 700216
rect 24302 700204 24308 700216
rect 24360 700204 24366 700256
rect 36722 700204 36728 700256
rect 36780 700244 36786 700256
rect 40494 700244 40500 700256
rect 36780 700216 40500 700244
rect 36780 700204 36786 700216
rect 40494 700204 40500 700216
rect 40552 700204 40558 700256
rect 69382 700204 69388 700256
rect 69440 700244 69446 700256
rect 72970 700244 72976 700256
rect 69440 700216 72976 700244
rect 69440 700204 69446 700216
rect 72970 700204 72976 700216
rect 73028 700204 73034 700256
rect 85758 700204 85764 700256
rect 85816 700244 85822 700256
rect 89162 700244 89168 700256
rect 85816 700216 89168 700244
rect 85816 700204 85822 700216
rect 89162 700204 89168 700216
rect 89220 700204 89226 700256
rect 134702 700204 134708 700256
rect 134760 700244 134766 700256
rect 137830 700244 137836 700256
rect 134760 700216 137836 700244
rect 134760 700204 134766 700216
rect 137830 700204 137836 700216
rect 137888 700204 137894 700256
rect 167362 700204 167368 700256
rect 167420 700244 167426 700256
rect 170306 700244 170312 700256
rect 167420 700216 170312 700244
rect 167420 700204 167426 700216
rect 170306 700204 170312 700216
rect 170364 700204 170370 700256
rect 183738 700204 183744 700256
rect 183796 700244 183802 700256
rect 186498 700244 186504 700256
rect 183796 700216 186504 700244
rect 183796 700204 183802 700216
rect 186498 700204 186504 700216
rect 186556 700204 186562 700256
rect 232774 700204 232780 700256
rect 232832 700244 232838 700256
rect 235166 700244 235172 700256
rect 232832 700216 235172 700244
rect 232832 700204 232838 700216
rect 235166 700204 235172 700216
rect 235224 700204 235230 700256
rect 249058 700204 249064 700256
rect 249116 700244 249122 700256
rect 251450 700244 251456 700256
rect 249116 700216 251456 700244
rect 249116 700204 249122 700216
rect 251450 700204 251456 700216
rect 251508 700204 251514 700256
rect 265434 700204 265440 700256
rect 265492 700244 265498 700256
rect 267642 700244 267648 700256
rect 265492 700216 267648 700244
rect 265492 700204 265498 700216
rect 267642 700204 267648 700216
rect 267700 700204 267706 700256
rect 281810 700204 281816 700256
rect 281868 700244 281874 700256
rect 283834 700244 283840 700256
rect 281868 700216 283840 700244
rect 281868 700204 281874 700216
rect 283834 700204 283840 700216
rect 283892 700204 283898 700256
rect 330754 700204 330760 700256
rect 330812 700244 330818 700256
rect 332502 700244 332508 700256
rect 330812 700216 332508 700244
rect 330812 700204 330818 700216
rect 332502 700204 332508 700216
rect 332560 700204 332566 700256
rect 347130 700204 347136 700256
rect 347188 700244 347194 700256
rect 348786 700244 348792 700256
rect 347188 700216 348792 700244
rect 347188 700204 347194 700216
rect 348786 700204 348792 700216
rect 348844 700204 348850 700256
rect 396166 700204 396172 700256
rect 396224 700244 396230 700256
rect 397454 700244 397460 700256
rect 396224 700216 397460 700244
rect 396224 700204 396230 700216
rect 397454 700204 397460 700216
rect 397512 700204 397518 700256
rect 428826 700204 428832 700256
rect 428884 700244 428890 700256
rect 429838 700244 429844 700256
rect 428884 700216 429844 700244
rect 428884 700204 428890 700216
rect 429838 700204 429844 700216
rect 429896 700204 429902 700256
rect 445202 700204 445208 700256
rect 445260 700244 445266 700256
rect 446122 700244 446128 700256
rect 445260 700216 446128 700244
rect 445260 700204 445266 700216
rect 446122 700204 446128 700216
rect 446180 700204 446186 700256
rect 461486 700204 461492 700256
rect 461544 700244 461550 700256
rect 462314 700244 462320 700256
rect 461544 700216 462320 700244
rect 461544 700204 461550 700216
rect 462314 700204 462320 700216
rect 462372 700204 462378 700256
rect 118418 700136 118424 700188
rect 118476 700176 118482 700188
rect 121638 700176 121644 700188
rect 118476 700148 121644 700176
rect 118476 700136 118482 700148
rect 121638 700136 121644 700148
rect 121696 700136 121702 700188
rect 216398 700136 216404 700188
rect 216456 700176 216462 700188
rect 218974 700176 218980 700188
rect 216456 700148 218980 700176
rect 216456 700136 216462 700148
rect 218974 700136 218980 700148
rect 219032 700136 219038 700188
rect 298002 700136 298008 700188
rect 298060 700176 298066 700188
rect 300118 700176 300124 700188
rect 298060 700148 300124 700176
rect 298060 700136 298066 700148
rect 300118 700136 300124 700148
rect 300176 700136 300182 700188
rect 477862 700136 477868 700188
rect 477920 700176 477926 700188
rect 478506 700176 478512 700188
rect 477920 700148 478512 700176
rect 477920 700136 477926 700148
rect 478506 700136 478512 700148
rect 478564 700136 478570 700188
rect 494238 700136 494244 700188
rect 494296 700176 494302 700188
rect 494790 700176 494796 700188
rect 494296 700148 494796 700176
rect 494296 700136 494302 700148
rect 494790 700136 494796 700148
rect 494848 700136 494854 700188
rect 379790 699864 379796 699916
rect 379848 699904 379854 699916
rect 381170 699904 381176 699916
rect 379848 699876 381176 699904
rect 379848 699864 379854 699876
rect 381170 699864 381176 699876
rect 381228 699864 381234 699916
rect 576762 698232 576768 698284
rect 576820 698272 576826 698284
rect 580166 698272 580172 698284
rect 576820 698244 580172 698272
rect 576820 698232 576826 698244
rect 580166 698232 580172 698244
rect 580224 698232 580230 698284
rect 4014 698164 4020 698216
rect 4072 698204 4078 698216
rect 8110 698204 8116 698216
rect 4072 698176 8116 698204
rect 4072 698164 4078 698176
rect 8110 698164 8116 698176
rect 8168 698164 8174 698216
rect 578326 644512 578332 644564
rect 578384 644552 578390 644564
rect 580902 644552 580908 644564
rect 578384 644524 580908 644552
rect 578384 644512 578390 644524
rect 580902 644512 580908 644524
rect 580960 644512 580966 644564
rect 578878 257796 578884 257848
rect 578936 257836 578942 257848
rect 580902 257836 580908 257848
rect 578936 257808 580908 257836
rect 578936 257796 578942 257808
rect 580902 257796 580908 257808
rect 580960 257796 580966 257848
rect 578510 151444 578516 151496
rect 578568 151484 578574 151496
rect 580902 151484 580908 151496
rect 578568 151456 580908 151484
rect 578568 151444 578574 151456
rect 580902 151444 580908 151456
rect 580960 151444 580966 151496
rect 578326 44956 578332 45008
rect 578384 44996 578390 45008
rect 579982 44996 579988 45008
rect 578384 44968 579988 44996
rect 578384 44956 578390 44968
rect 579982 44956 579988 44968
rect 580040 44956 580046 45008
rect 576854 5516 576860 5568
rect 576912 5556 576918 5568
rect 579614 5556 579620 5568
rect 576912 5528 579620 5556
rect 576912 5516 576918 5528
rect 579614 5516 579620 5528
rect 579672 5516 579678 5568
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 14502 3924 14508 3936
rect 11204 3896 14508 3924
rect 11204 3884 11210 3896
rect 14502 3884 14508 3896
rect 14560 3884 14566 3936
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 17998 3924 18004 3936
rect 14792 3896 18004 3924
rect 14792 3884 14798 3896
rect 17998 3884 18004 3896
rect 18056 3884 18062 3936
rect 20622 3884 20628 3936
rect 20680 3924 20686 3936
rect 23794 3924 23800 3936
rect 20680 3896 23800 3924
rect 20680 3884 20686 3896
rect 23794 3884 23800 3896
rect 23852 3884 23858 3936
rect 24210 3884 24216 3936
rect 24268 3924 24274 3936
rect 27290 3924 27296 3936
rect 24268 3896 27296 3924
rect 24268 3884 24274 3896
rect 27290 3884 27296 3896
rect 27348 3884 27354 3936
rect 27706 3884 27712 3936
rect 27764 3924 27770 3936
rect 30694 3924 30700 3936
rect 27764 3896 30700 3924
rect 27764 3884 27770 3896
rect 30694 3884 30700 3896
rect 30752 3884 30758 3936
rect 32398 3884 32404 3936
rect 32456 3924 32462 3936
rect 35386 3924 35392 3936
rect 32456 3896 35392 3924
rect 32456 3884 32462 3896
rect 35386 3884 35392 3896
rect 35444 3884 35450 3936
rect 38378 3884 38384 3936
rect 38436 3924 38442 3936
rect 41182 3924 41188 3936
rect 38436 3896 41188 3924
rect 38436 3884 38442 3896
rect 41182 3884 41188 3896
rect 41240 3884 41246 3936
rect 43070 3884 43076 3936
rect 43128 3924 43134 3936
rect 45782 3924 45788 3936
rect 43128 3896 45788 3924
rect 43128 3884 43134 3896
rect 45782 3884 45788 3896
rect 45840 3884 45846 3936
rect 46658 3884 46664 3936
rect 46716 3924 46722 3936
rect 49278 3924 49284 3936
rect 46716 3896 49284 3924
rect 46716 3884 46722 3896
rect 49278 3884 49284 3896
rect 49336 3884 49342 3936
rect 50154 3884 50160 3936
rect 50212 3924 50218 3936
rect 52774 3924 52780 3936
rect 50212 3896 52780 3924
rect 50212 3884 50218 3896
rect 52774 3884 52780 3896
rect 52832 3884 52838 3936
rect 56042 3884 56048 3936
rect 56100 3924 56106 3936
rect 58570 3924 58576 3936
rect 56100 3896 58576 3924
rect 56100 3884 56106 3896
rect 58570 3884 58576 3896
rect 58628 3884 58634 3936
rect 72602 3884 72608 3936
rect 72660 3924 72666 3936
rect 74854 3924 74860 3936
rect 72660 3896 74860 3924
rect 72660 3884 72666 3896
rect 74854 3884 74860 3896
rect 74912 3884 74918 3936
rect 247630 3884 247636 3936
rect 247688 3924 247694 3936
rect 248598 3924 248604 3936
rect 247688 3896 248604 3924
rect 247688 3884 247694 3896
rect 248598 3884 248604 3896
rect 248656 3884 248662 3936
rect 285902 3884 285908 3936
rect 285960 3924 285966 3936
rect 287790 3924 287796 3936
rect 285960 3896 287796 3924
rect 285960 3884 285966 3896
rect 287790 3884 287796 3896
rect 287848 3884 287854 3936
rect 1670 3816 1676 3868
rect 1728 3856 1734 3868
rect 5210 3856 5216 3868
rect 1728 3828 5216 3856
rect 1728 3816 1734 3828
rect 5210 3816 5216 3828
rect 5268 3816 5274 3868
rect 13538 3816 13544 3868
rect 13596 3856 13602 3868
rect 16802 3856 16808 3868
rect 13596 3828 16808 3856
rect 13596 3816 13602 3828
rect 16802 3816 16808 3828
rect 16860 3816 16866 3868
rect 19426 3816 19432 3868
rect 19484 3856 19490 3868
rect 22598 3856 22604 3868
rect 19484 3828 22604 3856
rect 19484 3816 19490 3828
rect 22598 3816 22604 3828
rect 22656 3816 22662 3868
rect 23014 3816 23020 3868
rect 23072 3856 23078 3868
rect 26094 3856 26100 3868
rect 23072 3828 26100 3856
rect 23072 3816 23078 3828
rect 26094 3816 26100 3828
rect 26152 3816 26158 3868
rect 26510 3816 26516 3868
rect 26568 3856 26574 3868
rect 29590 3856 29596 3868
rect 26568 3828 29596 3856
rect 26568 3816 26574 3828
rect 29590 3816 29596 3828
rect 29648 3816 29654 3868
rect 30098 3816 30104 3868
rect 30156 3856 30162 3868
rect 33086 3856 33092 3868
rect 30156 3828 33092 3856
rect 30156 3816 30162 3828
rect 33086 3816 33092 3828
rect 33144 3816 33150 3868
rect 33594 3816 33600 3868
rect 33652 3856 33658 3868
rect 36582 3856 36588 3868
rect 33652 3828 36588 3856
rect 33652 3816 33658 3828
rect 36582 3816 36588 3828
rect 36640 3816 36646 3868
rect 37182 3816 37188 3868
rect 37240 3856 37246 3868
rect 39986 3856 39992 3868
rect 37240 3828 39992 3856
rect 37240 3816 37246 3828
rect 39986 3816 39992 3828
rect 40044 3816 40050 3868
rect 41874 3816 41880 3868
rect 41932 3856 41938 3868
rect 44678 3856 44684 3868
rect 41932 3828 44684 3856
rect 41932 3816 41938 3828
rect 44678 3816 44684 3828
rect 44736 3816 44742 3868
rect 45462 3816 45468 3868
rect 45520 3856 45526 3868
rect 48174 3856 48180 3868
rect 45520 3828 48180 3856
rect 45520 3816 45526 3828
rect 48174 3816 48180 3828
rect 48232 3816 48238 3868
rect 48958 3816 48964 3868
rect 49016 3856 49022 3868
rect 51578 3856 51584 3868
rect 49016 3828 51584 3856
rect 49016 3816 49022 3828
rect 51578 3816 51584 3828
rect 51636 3816 51642 3868
rect 53742 3816 53748 3868
rect 53800 3856 53806 3868
rect 56270 3856 56276 3868
rect 53800 3828 56276 3856
rect 53800 3816 53806 3828
rect 56270 3816 56276 3828
rect 56328 3816 56334 3868
rect 57238 3816 57244 3868
rect 57296 3856 57302 3868
rect 59766 3856 59772 3868
rect 57296 3828 59772 3856
rect 57296 3816 57302 3828
rect 59766 3816 59772 3828
rect 59824 3816 59830 3868
rect 71498 3816 71504 3868
rect 71556 3856 71562 3868
rect 73658 3856 73664 3868
rect 71556 3828 73664 3856
rect 71556 3816 71562 3828
rect 73658 3816 73664 3828
rect 73716 3816 73722 3868
rect 78582 3816 78588 3868
rect 78640 3856 78646 3868
rect 80650 3856 80656 3868
rect 78640 3828 80656 3856
rect 78640 3816 78646 3828
rect 80650 3816 80656 3828
rect 80708 3816 80714 3868
rect 80882 3816 80888 3868
rect 80940 3856 80946 3868
rect 82950 3856 82956 3868
rect 80940 3828 82956 3856
rect 80940 3816 80946 3828
rect 82950 3816 82956 3828
rect 83008 3816 83014 3868
rect 87966 3816 87972 3868
rect 88024 3856 88030 3868
rect 89942 3856 89948 3868
rect 88024 3828 89948 3856
rect 88024 3816 88030 3828
rect 89942 3816 89948 3828
rect 90000 3816 90006 3868
rect 96246 3816 96252 3868
rect 96304 3856 96310 3868
rect 98038 3856 98044 3868
rect 96304 3828 98044 3856
rect 96304 3816 96310 3828
rect 98038 3816 98044 3828
rect 98096 3816 98102 3868
rect 244134 3816 244140 3868
rect 244192 3856 244198 3868
rect 245194 3856 245200 3868
rect 244192 3828 245200 3856
rect 244192 3816 244198 3828
rect 245194 3816 245200 3828
rect 245252 3816 245258 3868
rect 256922 3816 256928 3868
rect 256980 3856 256986 3868
rect 258258 3856 258264 3868
rect 256980 3828 258264 3856
rect 256980 3816 256986 3828
rect 258258 3816 258264 3828
rect 258316 3816 258322 3868
rect 259222 3816 259228 3868
rect 259280 3856 259286 3868
rect 260650 3856 260656 3868
rect 259280 3828 260656 3856
rect 259280 3816 259286 3828
rect 260650 3816 260656 3828
rect 260708 3816 260714 3868
rect 261614 3816 261620 3868
rect 261672 3856 261678 3868
rect 262950 3856 262956 3868
rect 261672 3828 262956 3856
rect 261672 3816 261678 3828
rect 262950 3816 262956 3828
rect 263008 3816 263014 3868
rect 263914 3816 263920 3868
rect 263972 3856 263978 3868
rect 265342 3856 265348 3868
rect 263972 3828 265348 3856
rect 263972 3816 263978 3828
rect 265342 3816 265348 3828
rect 265400 3816 265406 3868
rect 268514 3816 268520 3868
rect 268572 3856 268578 3868
rect 270034 3856 270040 3868
rect 268572 3828 270040 3856
rect 268572 3816 268578 3828
rect 270034 3816 270040 3828
rect 270092 3816 270098 3868
rect 270814 3816 270820 3868
rect 270872 3856 270878 3868
rect 272426 3856 272432 3868
rect 270872 3828 272432 3856
rect 270872 3816 270878 3828
rect 272426 3816 272432 3828
rect 272484 3816 272490 3868
rect 275506 3816 275512 3868
rect 275564 3856 275570 3868
rect 277118 3856 277124 3868
rect 275564 3828 277124 3856
rect 275564 3816 275570 3828
rect 277118 3816 277124 3828
rect 277176 3816 277182 3868
rect 277806 3816 277812 3868
rect 277864 3856 277870 3868
rect 279510 3856 279516 3868
rect 277864 3828 279516 3856
rect 277864 3816 277870 3828
rect 279510 3816 279516 3828
rect 279568 3816 279574 3868
rect 284798 3816 284804 3868
rect 284856 3856 284862 3868
rect 286594 3856 286600 3868
rect 284856 3828 286600 3856
rect 284856 3816 284862 3828
rect 286594 3816 286600 3828
rect 286652 3816 286658 3868
rect 292894 3816 292900 3868
rect 292952 3856 292958 3868
rect 294874 3856 294880 3868
rect 292952 3828 294880 3856
rect 292952 3816 292958 3828
rect 294874 3816 294880 3828
rect 294932 3816 294938 3868
rect 299886 3816 299892 3868
rect 299944 3856 299950 3868
rect 301958 3856 301964 3868
rect 299944 3828 301964 3856
rect 299944 3816 299950 3828
rect 301958 3816 301964 3828
rect 302016 3816 302022 3868
rect 306786 3816 306792 3868
rect 306844 3856 306850 3868
rect 309042 3856 309048 3868
rect 306844 3828 309048 3856
rect 306844 3816 306850 3828
rect 309042 3816 309048 3828
rect 309100 3816 309106 3868
rect 566 3748 572 3800
rect 624 3788 630 3800
rect 4106 3788 4112 3800
rect 624 3760 4112 3788
rect 624 3748 630 3760
rect 4106 3748 4112 3760
rect 4164 3748 4170 3800
rect 7650 3748 7656 3800
rect 7708 3788 7714 3800
rect 11006 3788 11012 3800
rect 7708 3760 11012 3788
rect 7708 3748 7714 3760
rect 11006 3748 11012 3760
rect 11064 3748 11070 3800
rect 12342 3748 12348 3800
rect 12400 3788 12406 3800
rect 15698 3788 15704 3800
rect 12400 3760 15704 3788
rect 12400 3748 12406 3760
rect 15698 3748 15704 3760
rect 15756 3748 15762 3800
rect 15930 3748 15936 3800
rect 15988 3788 15994 3800
rect 19102 3788 19108 3800
rect 15988 3760 19108 3788
rect 15988 3748 15994 3760
rect 19102 3748 19108 3760
rect 19160 3748 19166 3800
rect 21818 3748 21824 3800
rect 21876 3788 21882 3800
rect 24898 3788 24904 3800
rect 21876 3760 24904 3788
rect 21876 3748 21882 3760
rect 24898 3748 24904 3760
rect 24956 3748 24962 3800
rect 25314 3748 25320 3800
rect 25372 3788 25378 3800
rect 28394 3788 28400 3800
rect 25372 3760 28400 3788
rect 25372 3748 25378 3760
rect 28394 3748 28400 3760
rect 28452 3748 28458 3800
rect 31294 3748 31300 3800
rect 31352 3788 31358 3800
rect 34190 3788 34196 3800
rect 31352 3760 34196 3788
rect 31352 3748 31358 3760
rect 34190 3748 34196 3760
rect 34248 3748 34254 3800
rect 34790 3748 34796 3800
rect 34848 3788 34854 3800
rect 37686 3788 37692 3800
rect 34848 3760 37692 3788
rect 34848 3748 34854 3760
rect 37686 3748 37692 3760
rect 37744 3748 37750 3800
rect 40678 3748 40684 3800
rect 40736 3788 40742 3800
rect 43482 3788 43488 3800
rect 40736 3760 43488 3788
rect 40736 3748 40742 3760
rect 43482 3748 43488 3760
rect 43540 3748 43546 3800
rect 44266 3748 44272 3800
rect 44324 3788 44330 3800
rect 46978 3788 46984 3800
rect 44324 3760 46984 3788
rect 44324 3748 44330 3760
rect 46978 3748 46984 3760
rect 47036 3748 47042 3800
rect 47854 3748 47860 3800
rect 47912 3788 47918 3800
rect 50474 3788 50480 3800
rect 47912 3760 50480 3788
rect 47912 3748 47918 3760
rect 50474 3748 50480 3760
rect 50532 3748 50538 3800
rect 51350 3748 51356 3800
rect 51408 3788 51414 3800
rect 53970 3788 53976 3800
rect 51408 3760 53976 3788
rect 51408 3748 51414 3760
rect 53970 3748 53976 3760
rect 54028 3748 54034 3800
rect 54938 3748 54944 3800
rect 54996 3788 55002 3800
rect 57374 3788 57380 3800
rect 54996 3760 57380 3788
rect 54996 3748 55002 3760
rect 57374 3748 57380 3760
rect 57432 3748 57438 3800
rect 58434 3748 58440 3800
rect 58492 3788 58498 3800
rect 60870 3788 60876 3800
rect 58492 3760 60876 3788
rect 58492 3748 58498 3760
rect 60870 3748 60876 3760
rect 60928 3748 60934 3800
rect 64322 3748 64328 3800
rect 64380 3788 64386 3800
rect 66666 3788 66672 3800
rect 64380 3760 66672 3788
rect 64380 3748 64386 3760
rect 66666 3748 66672 3760
rect 66724 3748 66730 3800
rect 67082 3748 67088 3800
rect 67140 3788 67146 3800
rect 69058 3788 69064 3800
rect 67140 3760 69064 3788
rect 67140 3748 67146 3760
rect 69058 3748 69064 3760
rect 69116 3748 69122 3800
rect 70302 3748 70308 3800
rect 70360 3788 70366 3800
rect 72462 3788 72468 3800
rect 70360 3760 72468 3788
rect 70360 3748 70366 3760
rect 72462 3748 72468 3760
rect 72520 3748 72526 3800
rect 73798 3748 73804 3800
rect 73856 3788 73862 3800
rect 75958 3788 75964 3800
rect 73856 3760 75964 3788
rect 73856 3748 73862 3760
rect 75958 3748 75964 3760
rect 76016 3748 76022 3800
rect 79686 3748 79692 3800
rect 79744 3788 79750 3800
rect 81754 3788 81760 3800
rect 79744 3760 81760 3788
rect 79744 3748 79750 3760
rect 81754 3748 81760 3760
rect 81812 3748 81818 3800
rect 86862 3748 86868 3800
rect 86920 3788 86926 3800
rect 88746 3788 88752 3800
rect 86920 3760 88752 3788
rect 86920 3748 86926 3760
rect 88746 3748 88752 3760
rect 88804 3748 88810 3800
rect 95142 3748 95148 3800
rect 95200 3788 95206 3800
rect 96842 3788 96848 3800
rect 95200 3760 96848 3788
rect 95200 3748 95206 3760
rect 96842 3748 96848 3760
rect 96900 3748 96906 3800
rect 103330 3748 103336 3800
rect 103388 3788 103394 3800
rect 104938 3788 104944 3800
rect 103388 3760 104944 3788
rect 103388 3748 103394 3760
rect 104938 3748 104944 3760
rect 104996 3748 105002 3800
rect 216350 3748 216356 3800
rect 216408 3788 216414 3800
rect 216858 3788 216864 3800
rect 216408 3760 216864 3788
rect 216408 3748 216414 3760
rect 216858 3748 216864 3760
rect 216916 3748 216922 3800
rect 222146 3748 222152 3800
rect 222204 3788 222210 3800
rect 222746 3788 222752 3800
rect 222204 3760 222752 3788
rect 222204 3748 222210 3760
rect 222746 3748 222752 3760
rect 222804 3748 222810 3800
rect 224446 3748 224452 3800
rect 224504 3788 224510 3800
rect 225138 3788 225144 3800
rect 224504 3760 225144 3788
rect 224504 3748 224510 3760
rect 225138 3748 225144 3760
rect 225196 3748 225202 3800
rect 230242 3748 230248 3800
rect 230300 3788 230306 3800
rect 231026 3788 231032 3800
rect 230300 3760 231032 3788
rect 230300 3748 230306 3760
rect 231026 3748 231032 3760
rect 231084 3748 231090 3800
rect 231438 3748 231444 3800
rect 231496 3788 231502 3800
rect 232222 3788 232228 3800
rect 231496 3760 232228 3788
rect 231496 3748 231502 3760
rect 232222 3748 232228 3760
rect 232280 3748 232286 3800
rect 232542 3748 232548 3800
rect 232600 3788 232606 3800
rect 233418 3788 233424 3800
rect 232600 3760 233424 3788
rect 232600 3748 232606 3760
rect 233418 3748 233424 3760
rect 233476 3748 233482 3800
rect 233738 3748 233744 3800
rect 233796 3788 233802 3800
rect 234614 3788 234620 3800
rect 233796 3760 234620 3788
rect 233796 3748 233802 3760
rect 234614 3748 234620 3760
rect 234672 3748 234678 3800
rect 237234 3748 237240 3800
rect 237292 3788 237298 3800
rect 238110 3788 238116 3800
rect 237292 3760 238116 3788
rect 237292 3748 237298 3760
rect 238110 3748 238116 3760
rect 238168 3748 238174 3800
rect 238338 3748 238344 3800
rect 238396 3788 238402 3800
rect 239306 3788 239312 3800
rect 238396 3760 239312 3788
rect 238396 3748 238402 3760
rect 239306 3748 239312 3760
rect 239364 3748 239370 3800
rect 239534 3748 239540 3800
rect 239592 3788 239598 3800
rect 240502 3788 240508 3800
rect 239592 3760 240508 3788
rect 239592 3748 239598 3760
rect 240502 3748 240508 3760
rect 240560 3748 240566 3800
rect 240730 3748 240736 3800
rect 240788 3788 240794 3800
rect 241698 3788 241704 3800
rect 240788 3760 241704 3788
rect 240788 3748 240794 3760
rect 241698 3748 241704 3760
rect 241756 3748 241762 3800
rect 241834 3748 241840 3800
rect 241892 3788 241898 3800
rect 242894 3788 242900 3800
rect 241892 3760 242900 3788
rect 241892 3748 241898 3760
rect 242894 3748 242900 3760
rect 242952 3748 242958 3800
rect 245330 3748 245336 3800
rect 245388 3788 245394 3800
rect 246390 3788 246396 3800
rect 245388 3760 246396 3788
rect 245388 3748 245394 3760
rect 246390 3748 246396 3760
rect 246448 3748 246454 3800
rect 246526 3748 246532 3800
rect 246584 3788 246590 3800
rect 247586 3788 247592 3800
rect 246584 3760 247592 3788
rect 246584 3748 246590 3760
rect 247586 3748 247592 3760
rect 247644 3748 247650 3800
rect 250022 3748 250028 3800
rect 250080 3788 250086 3800
rect 251174 3788 251180 3800
rect 250080 3760 251180 3788
rect 250080 3748 250086 3760
rect 251174 3748 251180 3760
rect 251232 3748 251238 3800
rect 252322 3748 252328 3800
rect 252380 3788 252386 3800
rect 253474 3788 253480 3800
rect 252380 3760 253480 3788
rect 252380 3748 252386 3760
rect 253474 3748 253480 3760
rect 253532 3748 253538 3800
rect 255818 3748 255824 3800
rect 255876 3788 255882 3800
rect 257062 3788 257068 3800
rect 255876 3760 257068 3788
rect 255876 3748 255882 3760
rect 257062 3748 257068 3760
rect 257120 3748 257126 3800
rect 258118 3748 258124 3800
rect 258176 3788 258182 3800
rect 259454 3788 259460 3800
rect 258176 3760 259460 3788
rect 258176 3748 258182 3760
rect 259454 3748 259460 3760
rect 259512 3748 259518 3800
rect 260418 3748 260424 3800
rect 260476 3788 260482 3800
rect 261754 3788 261760 3800
rect 260476 3760 261760 3788
rect 260476 3748 260482 3760
rect 261754 3748 261760 3760
rect 261812 3748 261818 3800
rect 262718 3748 262724 3800
rect 262776 3788 262782 3800
rect 264146 3788 264152 3800
rect 262776 3760 264152 3788
rect 262776 3748 262782 3760
rect 264146 3748 264152 3760
rect 264204 3748 264210 3800
rect 265018 3748 265024 3800
rect 265076 3788 265082 3800
rect 266538 3788 266544 3800
rect 265076 3760 266544 3788
rect 265076 3748 265082 3760
rect 266538 3748 266544 3760
rect 266596 3748 266602 3800
rect 267410 3748 267416 3800
rect 267468 3788 267474 3800
rect 268838 3788 268844 3800
rect 267468 3760 268844 3788
rect 267468 3748 267474 3760
rect 268838 3748 268844 3760
rect 268896 3748 268902 3800
rect 269710 3748 269716 3800
rect 269768 3788 269774 3800
rect 271230 3788 271236 3800
rect 269768 3760 271236 3788
rect 269768 3748 269774 3760
rect 271230 3748 271236 3760
rect 271288 3748 271294 3800
rect 272010 3748 272016 3800
rect 272068 3788 272074 3800
rect 273622 3788 273628 3800
rect 272068 3760 273628 3788
rect 272068 3748 272074 3760
rect 273622 3748 273628 3760
rect 273680 3748 273686 3800
rect 276702 3748 276708 3800
rect 276760 3788 276766 3800
rect 278314 3788 278320 3800
rect 276760 3760 278320 3788
rect 276760 3748 276766 3760
rect 278314 3748 278320 3760
rect 278372 3748 278378 3800
rect 279002 3748 279008 3800
rect 279060 3788 279066 3800
rect 280706 3788 280712 3800
rect 279060 3760 280712 3788
rect 279060 3748 279066 3760
rect 280706 3748 280712 3760
rect 280764 3748 280770 3800
rect 283602 3748 283608 3800
rect 283660 3788 283666 3800
rect 285398 3788 285404 3800
rect 283660 3760 285404 3788
rect 283660 3748 283666 3760
rect 285398 3748 285404 3760
rect 285456 3748 285462 3800
rect 287098 3748 287104 3800
rect 287156 3788 287162 3800
rect 288986 3788 288992 3800
rect 287156 3760 288992 3788
rect 287156 3748 287162 3760
rect 288986 3748 288992 3760
rect 289044 3748 289050 3800
rect 291698 3748 291704 3800
rect 291756 3788 291762 3800
rect 293678 3788 293684 3800
rect 291756 3760 293684 3788
rect 291756 3748 291762 3760
rect 293678 3748 293684 3760
rect 293736 3748 293742 3800
rect 294090 3748 294096 3800
rect 294148 3788 294154 3800
rect 296070 3788 296076 3800
rect 294148 3760 296076 3788
rect 294148 3748 294154 3760
rect 296070 3748 296076 3760
rect 296128 3748 296134 3800
rect 298690 3748 298696 3800
rect 298748 3788 298754 3800
rect 300762 3788 300768 3800
rect 298748 3760 300768 3788
rect 298748 3748 298754 3760
rect 300762 3748 300768 3760
rect 300820 3748 300826 3800
rect 300990 3748 300996 3800
rect 301048 3788 301054 3800
rect 303154 3788 303160 3800
rect 301048 3760 303160 3788
rect 301048 3748 301054 3760
rect 303154 3748 303160 3760
rect 303212 3748 303218 3800
rect 307982 3748 307988 3800
rect 308040 3788 308046 3800
rect 310238 3788 310244 3800
rect 308040 3760 310244 3788
rect 308040 3748 308046 3760
rect 310238 3748 310244 3760
rect 310296 3748 310302 3800
rect 316078 3748 316084 3800
rect 316136 3788 316142 3800
rect 318518 3788 318524 3800
rect 316136 3760 318524 3788
rect 316136 3748 316142 3760
rect 318518 3748 318524 3760
rect 318576 3748 318582 3800
rect 323070 3748 323076 3800
rect 323128 3788 323134 3800
rect 325602 3788 325608 3800
rect 323128 3760 325608 3788
rect 323128 3748 323134 3760
rect 325602 3748 325608 3760
rect 325660 3748 325666 3800
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 9858 3040 9864 3052
rect 6512 3012 9864 3040
rect 6512 3000 6518 3012
rect 9858 3000 9864 3012
rect 9916 3000 9922 3052
rect 63218 3000 63224 3052
rect 63276 3040 63282 3052
rect 65518 3040 65524 3052
rect 63276 3012 65524 3040
rect 63276 3000 63282 3012
rect 65518 3000 65524 3012
rect 65576 3000 65582 3052
rect 18230 2864 18236 2916
rect 18288 2904 18294 2916
rect 21450 2904 21456 2916
rect 18288 2876 21456 2904
rect 18288 2864 18294 2876
rect 21450 2864 21456 2876
rect 21508 2864 21514 2916
rect 253382 2864 253388 2916
rect 253440 2904 253446 2916
rect 254670 2904 254676 2916
rect 253440 2876 254676 2904
rect 253440 2864 253446 2876
rect 254670 2864 254676 2876
rect 254728 2864 254734 2916
rect 4062 2796 4068 2848
rect 4120 2836 4126 2848
rect 7466 2836 7472 2848
rect 4120 2808 7472 2836
rect 4120 2796 4126 2808
rect 7466 2796 7472 2808
rect 7524 2796 7530 2848
rect 9950 2796 9956 2848
rect 10008 2836 10014 2848
rect 13262 2836 13268 2848
rect 10008 2808 13268 2836
rect 10008 2796 10014 2808
rect 13262 2796 13268 2808
rect 13320 2796 13326 2848
rect 17034 2796 17040 2848
rect 17092 2836 17098 2848
rect 20254 2836 20260 2848
rect 17092 2808 20260 2836
rect 17092 2796 17098 2808
rect 20254 2796 20260 2808
rect 20312 2796 20318 2848
rect 28902 2796 28908 2848
rect 28960 2836 28966 2848
rect 31846 2836 31852 2848
rect 28960 2808 31852 2836
rect 28960 2796 28966 2808
rect 31846 2796 31852 2808
rect 31904 2796 31910 2848
rect 35986 2796 35992 2848
rect 36044 2836 36050 2848
rect 38838 2836 38844 2848
rect 36044 2808 38844 2836
rect 36044 2796 36050 2808
rect 38838 2796 38844 2808
rect 38896 2796 38902 2848
rect 39574 2796 39580 2848
rect 39632 2836 39638 2848
rect 42334 2836 42340 2848
rect 39632 2808 42340 2836
rect 39632 2796 39638 2808
rect 42334 2796 42340 2808
rect 42392 2796 42398 2848
rect 62022 2796 62028 2848
rect 62080 2836 62086 2848
rect 64414 2836 64420 2848
rect 62080 2808 64420 2836
rect 62080 2796 62086 2808
rect 64414 2796 64420 2808
rect 64472 2796 64478 2848
rect 65518 2796 65524 2848
rect 65576 2836 65582 2848
rect 67818 2836 67824 2848
rect 65576 2808 67824 2836
rect 65576 2796 65582 2808
rect 67818 2796 67824 2808
rect 67876 2796 67882 2848
rect 248874 2796 248880 2848
rect 248932 2836 248938 2848
rect 249978 2836 249984 2848
rect 248932 2808 249984 2836
rect 248932 2796 248938 2808
rect 249978 2796 249984 2808
rect 250036 2796 250042 2848
rect 251082 2796 251088 2848
rect 251140 2836 251146 2848
rect 252370 2836 252376 2848
rect 251140 2808 252376 2836
rect 251140 2796 251146 2808
rect 252370 2796 252376 2808
rect 252428 2796 252434 2848
rect 254578 2796 254584 2848
rect 254636 2836 254642 2848
rect 255866 2836 255872 2848
rect 254636 2808 255872 2836
rect 254636 2796 254642 2808
rect 255866 2796 255872 2808
rect 255924 2796 255930 2848
rect 309226 2796 309232 2848
rect 309284 2836 309290 2848
rect 311434 2836 311440 2848
rect 309284 2808 311440 2836
rect 309284 2796 309290 2808
rect 311434 2796 311440 2808
rect 311492 2796 311498 2848
rect 315022 2796 315028 2848
rect 315080 2836 315086 2848
rect 317322 2836 317328 2848
rect 315080 2808 317328 2836
rect 315080 2796 315086 2808
rect 317322 2796 317328 2808
rect 317380 2796 317386 2848
rect 411162 2796 411168 2848
rect 411220 2836 411226 2848
rect 415486 2836 415492 2848
rect 411220 2808 415492 2836
rect 411220 2796 411226 2808
rect 415486 2796 415492 2808
rect 415544 2796 415550 2848
rect 440142 2796 440148 2848
rect 440200 2836 440206 2848
rect 445018 2836 445024 2848
rect 440200 2808 445024 2836
rect 440200 2796 440206 2808
rect 445018 2796 445024 2808
rect 445076 2796 445082 2848
rect 449526 2796 449532 2848
rect 449584 2836 449590 2848
rect 454494 2836 454500 2848
rect 449584 2808 454500 2836
rect 449584 2796 449590 2808
rect 454494 2796 454500 2808
rect 454552 2796 454558 2848
rect 478506 2796 478512 2848
rect 478564 2836 478570 2848
rect 484026 2836 484032 2848
rect 478564 2808 484032 2836
rect 478564 2796 478570 2808
rect 484026 2796 484032 2808
rect 484084 2796 484090 2848
rect 3234 1300 3240 1352
rect 3292 1340 3298 1352
rect 6362 1340 6368 1352
rect 3292 1312 6368 1340
rect 3292 1300 3298 1312
rect 6362 1300 6368 1312
rect 6420 1300 6426 1352
rect 60826 1300 60832 1352
rect 60884 1340 60890 1352
rect 63310 1340 63316 1352
rect 60884 1312 63316 1340
rect 60884 1300 60890 1312
rect 63310 1300 63316 1312
rect 63368 1300 63374 1352
rect 67910 1300 67916 1352
rect 67968 1340 67974 1352
rect 70118 1340 70124 1352
rect 67968 1312 70124 1340
rect 67968 1300 67974 1312
rect 70118 1300 70124 1312
rect 70176 1300 70182 1352
rect 76190 1300 76196 1352
rect 76248 1340 76254 1352
rect 78214 1340 78220 1352
rect 76248 1312 78220 1340
rect 76248 1300 76254 1312
rect 78214 1300 78220 1312
rect 78272 1300 78278 1352
rect 83274 1300 83280 1352
rect 83332 1340 83338 1352
rect 85206 1340 85212 1352
rect 83332 1312 85212 1340
rect 83332 1300 83338 1312
rect 85206 1300 85212 1312
rect 85264 1300 85270 1352
rect 85666 1300 85672 1352
rect 85724 1340 85730 1352
rect 87506 1340 87512 1352
rect 85724 1312 87512 1340
rect 85724 1300 85730 1312
rect 87506 1300 87512 1312
rect 87564 1300 87570 1352
rect 89162 1300 89168 1352
rect 89220 1340 89226 1352
rect 91002 1340 91008 1352
rect 89220 1312 91008 1340
rect 89220 1300 89226 1312
rect 91002 1300 91008 1312
rect 91060 1300 91066 1352
rect 91554 1300 91560 1352
rect 91612 1340 91618 1352
rect 93302 1340 93308 1352
rect 91612 1312 93308 1340
rect 91612 1300 91618 1312
rect 93302 1300 93308 1312
rect 93360 1300 93366 1352
rect 93946 1300 93952 1352
rect 94004 1340 94010 1352
rect 95694 1340 95700 1352
rect 94004 1312 95700 1340
rect 94004 1300 94010 1312
rect 95694 1300 95700 1312
rect 95752 1300 95758 1352
rect 97442 1300 97448 1352
rect 97500 1340 97506 1352
rect 99098 1340 99104 1352
rect 97500 1312 99104 1340
rect 97500 1300 97506 1312
rect 99098 1300 99104 1312
rect 99156 1300 99162 1352
rect 101030 1300 101036 1352
rect 101088 1340 101094 1352
rect 102594 1340 102600 1352
rect 101088 1312 102600 1340
rect 101088 1300 101094 1312
rect 102594 1300 102600 1312
rect 102652 1300 102658 1352
rect 104526 1300 104532 1352
rect 104584 1340 104590 1352
rect 106090 1340 106096 1352
rect 104584 1312 106096 1340
rect 104584 1300 104590 1312
rect 106090 1300 106096 1312
rect 106148 1300 106154 1352
rect 106918 1300 106924 1352
rect 106976 1340 106982 1352
rect 108390 1340 108396 1352
rect 106976 1312 108396 1340
rect 106976 1300 106982 1312
rect 108390 1300 108396 1312
rect 108448 1300 108454 1352
rect 109310 1300 109316 1352
rect 109368 1340 109374 1352
rect 110690 1340 110696 1352
rect 109368 1312 110696 1340
rect 109368 1300 109374 1312
rect 110690 1300 110696 1312
rect 110748 1300 110754 1352
rect 112806 1300 112812 1352
rect 112864 1340 112870 1352
rect 114186 1340 114192 1352
rect 112864 1312 114192 1340
rect 112864 1300 112870 1312
rect 114186 1300 114192 1312
rect 114244 1300 114250 1352
rect 116394 1300 116400 1352
rect 116452 1340 116458 1352
rect 117682 1340 117688 1352
rect 116452 1312 117688 1340
rect 116452 1300 116458 1312
rect 117682 1300 117688 1312
rect 117740 1300 117746 1352
rect 119890 1300 119896 1352
rect 119948 1340 119954 1352
rect 121178 1340 121184 1352
rect 119948 1312 121184 1340
rect 119948 1300 119954 1312
rect 121178 1300 121184 1312
rect 121236 1300 121242 1352
rect 125870 1300 125876 1352
rect 125928 1340 125934 1352
rect 126974 1340 126980 1352
rect 125928 1312 126980 1340
rect 125928 1300 125934 1312
rect 126974 1300 126980 1312
rect 127032 1300 127038 1352
rect 129366 1300 129372 1352
rect 129424 1340 129430 1352
rect 130470 1340 130476 1352
rect 129424 1312 130476 1340
rect 129424 1300 129430 1312
rect 130470 1300 130476 1312
rect 130528 1300 130534 1352
rect 130562 1300 130568 1352
rect 130620 1340 130626 1352
rect 131574 1340 131580 1352
rect 130620 1312 131580 1340
rect 130620 1300 130626 1312
rect 131574 1300 131580 1312
rect 131632 1300 131638 1352
rect 131758 1300 131764 1352
rect 131816 1340 131822 1352
rect 132770 1340 132776 1352
rect 131816 1312 132776 1340
rect 131816 1300 131822 1312
rect 132770 1300 132776 1312
rect 132828 1300 132834 1352
rect 132954 1300 132960 1352
rect 133012 1340 133018 1352
rect 133966 1340 133972 1352
rect 133012 1312 133972 1340
rect 133012 1300 133018 1312
rect 133966 1300 133972 1312
rect 134024 1300 134030 1352
rect 137646 1300 137652 1352
rect 137704 1340 137710 1352
rect 138566 1340 138572 1352
rect 137704 1312 138572 1340
rect 137704 1300 137710 1312
rect 138566 1300 138572 1312
rect 138624 1300 138630 1352
rect 144730 1300 144736 1352
rect 144788 1340 144794 1352
rect 145558 1340 145564 1352
rect 144788 1312 145564 1340
rect 144788 1300 144794 1312
rect 145558 1300 145564 1312
rect 145616 1300 145622 1352
rect 145926 1300 145932 1352
rect 145984 1340 145990 1352
rect 146662 1340 146668 1352
rect 145984 1312 146668 1340
rect 145984 1300 145990 1312
rect 146662 1300 146668 1312
rect 146720 1300 146726 1352
rect 148318 1300 148324 1352
rect 148376 1340 148382 1352
rect 149054 1340 149060 1352
rect 148376 1312 149060 1340
rect 148376 1300 148382 1312
rect 149054 1300 149060 1312
rect 149112 1300 149118 1352
rect 154206 1300 154212 1352
rect 154264 1340 154270 1352
rect 154850 1340 154856 1352
rect 154264 1312 154856 1340
rect 154264 1300 154270 1312
rect 154850 1300 154856 1312
rect 154908 1300 154914 1352
rect 162486 1300 162492 1352
rect 162544 1340 162550 1352
rect 162946 1340 162952 1352
rect 162544 1312 162952 1340
rect 162544 1300 162550 1312
rect 162946 1300 162952 1312
rect 163004 1300 163010 1352
rect 266262 1300 266268 1352
rect 266320 1340 266326 1352
rect 267734 1340 267740 1352
rect 266320 1312 267740 1340
rect 266320 1300 266326 1312
rect 267734 1300 267740 1312
rect 267792 1300 267798 1352
rect 273162 1300 273168 1352
rect 273220 1340 273226 1352
rect 274818 1340 274824 1352
rect 273220 1312 274824 1340
rect 273220 1300 273226 1312
rect 274818 1300 274824 1312
rect 274876 1300 274882 1352
rect 280062 1300 280068 1352
rect 280120 1340 280126 1352
rect 281902 1340 281908 1352
rect 280120 1312 281908 1340
rect 280120 1300 280126 1312
rect 281902 1300 281908 1312
rect 281960 1300 281966 1352
rect 282546 1300 282552 1352
rect 282604 1340 282610 1352
rect 284294 1340 284300 1352
rect 282604 1312 284300 1340
rect 282604 1300 282610 1312
rect 284294 1300 284300 1312
rect 284352 1300 284358 1352
rect 288342 1300 288348 1352
rect 288400 1340 288406 1352
rect 290182 1340 290188 1352
rect 288400 1312 290188 1340
rect 288400 1300 288406 1312
rect 290182 1300 290188 1312
rect 290240 1300 290246 1352
rect 295242 1300 295248 1352
rect 295300 1340 295306 1352
rect 297266 1340 297272 1352
rect 295300 1312 297272 1340
rect 295300 1300 295306 1312
rect 297266 1300 297272 1312
rect 297324 1300 297330 1352
rect 297542 1300 297548 1352
rect 297600 1340 297606 1352
rect 299658 1340 299664 1352
rect 297600 1312 299664 1340
rect 297600 1300 297606 1312
rect 299658 1300 299664 1312
rect 299716 1300 299722 1352
rect 302142 1300 302148 1352
rect 302200 1340 302206 1352
rect 304350 1340 304356 1352
rect 302200 1312 304356 1340
rect 302200 1300 302206 1312
rect 304350 1300 304356 1312
rect 304408 1300 304414 1352
rect 305730 1300 305736 1352
rect 305788 1340 305794 1352
rect 307938 1340 307944 1352
rect 305788 1312 307944 1340
rect 305788 1300 305794 1312
rect 307938 1300 307944 1312
rect 307996 1300 308002 1352
rect 310330 1300 310336 1352
rect 310388 1340 310394 1352
rect 312630 1340 312636 1352
rect 310388 1312 312636 1340
rect 310388 1300 310394 1312
rect 312630 1300 312636 1312
rect 312688 1300 312694 1352
rect 313826 1300 313832 1352
rect 313884 1340 313890 1352
rect 316218 1340 316224 1352
rect 313884 1312 316224 1340
rect 313884 1300 313890 1312
rect 316218 1300 316224 1312
rect 316276 1300 316282 1352
rect 317230 1300 317236 1352
rect 317288 1340 317294 1352
rect 319714 1340 319720 1352
rect 317288 1312 319720 1340
rect 317288 1300 317294 1312
rect 319714 1300 319720 1312
rect 319772 1300 319778 1352
rect 321922 1300 321928 1352
rect 321980 1340 321986 1352
rect 324406 1340 324412 1352
rect 321980 1312 324412 1340
rect 321980 1300 321986 1312
rect 324406 1300 324412 1312
rect 324464 1300 324470 1352
rect 325418 1300 325424 1352
rect 325476 1340 325482 1352
rect 327994 1340 328000 1352
rect 325476 1312 328000 1340
rect 325476 1300 325482 1312
rect 327994 1300 328000 1312
rect 328052 1300 328058 1352
rect 328914 1300 328920 1352
rect 328972 1340 328978 1352
rect 331582 1340 331588 1352
rect 328972 1312 331588 1340
rect 328972 1300 328978 1312
rect 331582 1300 331588 1312
rect 331640 1300 331646 1352
rect 332410 1300 332416 1352
rect 332468 1340 332474 1352
rect 335078 1340 335084 1352
rect 332468 1312 335084 1340
rect 332468 1300 332474 1312
rect 335078 1300 335084 1312
rect 335136 1300 335142 1352
rect 335906 1300 335912 1352
rect 335964 1340 335970 1352
rect 338666 1340 338672 1352
rect 335964 1312 338672 1340
rect 335964 1300 335970 1312
rect 338666 1300 338672 1312
rect 338724 1300 338730 1352
rect 339310 1300 339316 1352
rect 339368 1340 339374 1352
rect 342162 1340 342168 1352
rect 339368 1312 342168 1340
rect 339368 1300 339374 1312
rect 342162 1300 342168 1312
rect 342220 1300 342226 1352
rect 345106 1300 345112 1352
rect 345164 1340 345170 1352
rect 348050 1340 348056 1352
rect 345164 1312 348056 1340
rect 345164 1300 345170 1312
rect 348050 1300 348056 1312
rect 348108 1300 348114 1352
rect 349798 1300 349804 1352
rect 349856 1340 349862 1352
rect 352834 1340 352840 1352
rect 349856 1312 352840 1340
rect 349856 1300 349862 1312
rect 352834 1300 352840 1312
rect 352892 1300 352898 1352
rect 353202 1300 353208 1352
rect 353260 1340 353266 1352
rect 356330 1340 356336 1352
rect 353260 1312 356336 1340
rect 353260 1300 353266 1312
rect 356330 1300 356336 1312
rect 356388 1300 356394 1352
rect 356698 1300 356704 1352
rect 356756 1340 356762 1352
rect 359918 1340 359924 1352
rect 356756 1312 359924 1340
rect 356756 1300 356762 1312
rect 359918 1300 359924 1312
rect 359976 1300 359982 1352
rect 362586 1300 362592 1352
rect 362644 1340 362650 1352
rect 365806 1340 365812 1352
rect 362644 1312 365812 1340
rect 362644 1300 362650 1312
rect 365806 1300 365812 1312
rect 365864 1300 365870 1352
rect 367186 1300 367192 1352
rect 367244 1340 367250 1352
rect 370590 1340 370596 1352
rect 367244 1312 370596 1340
rect 367244 1300 367250 1312
rect 370590 1300 370596 1312
rect 370648 1300 370654 1352
rect 370682 1300 370688 1352
rect 370740 1340 370746 1352
rect 374086 1340 374092 1352
rect 370740 1312 374092 1340
rect 370740 1300 370746 1312
rect 374086 1300 374092 1312
rect 374144 1300 374150 1352
rect 376386 1300 376392 1352
rect 376444 1340 376450 1352
rect 379974 1340 379980 1352
rect 376444 1312 379980 1340
rect 376444 1300 376450 1312
rect 379974 1300 379980 1312
rect 380032 1300 380038 1352
rect 385770 1300 385776 1352
rect 385828 1340 385834 1352
rect 389450 1340 389456 1352
rect 385828 1312 389456 1340
rect 385828 1300 385834 1312
rect 389450 1300 389456 1312
rect 389508 1300 389514 1352
rect 395062 1300 395068 1352
rect 395120 1340 395126 1352
rect 398926 1340 398932 1352
rect 395120 1312 398932 1340
rect 395120 1300 395126 1312
rect 398926 1300 398932 1312
rect 398984 1300 398990 1352
rect 399662 1300 399668 1352
rect 399720 1340 399726 1352
rect 403618 1340 403624 1352
rect 399720 1312 403624 1340
rect 399720 1300 399726 1312
rect 403618 1300 403624 1312
rect 403676 1300 403682 1352
rect 405458 1300 405464 1352
rect 405516 1340 405522 1352
rect 409598 1340 409604 1352
rect 405516 1312 409604 1340
rect 405516 1300 405522 1312
rect 409598 1300 409604 1312
rect 409656 1300 409662 1352
rect 415946 1300 415952 1352
rect 416004 1340 416010 1352
rect 420178 1340 420184 1352
rect 416004 1312 420184 1340
rect 416004 1300 416010 1312
rect 420178 1300 420184 1312
rect 420236 1300 420242 1352
rect 427538 1300 427544 1352
rect 427596 1340 427602 1352
rect 431862 1340 431868 1352
rect 427596 1312 431868 1340
rect 427596 1300 427602 1312
rect 431862 1300 431868 1312
rect 431920 1300 431926 1352
rect 433242 1300 433248 1352
rect 433300 1340 433306 1352
rect 437842 1340 437848 1352
rect 433300 1312 437848 1340
rect 433300 1300 433306 1312
rect 437842 1300 437848 1312
rect 437900 1300 437906 1352
rect 442626 1300 442632 1352
rect 442684 1340 442690 1352
rect 447410 1340 447416 1352
rect 442684 1312 447416 1340
rect 442684 1300 442690 1312
rect 447410 1300 447416 1312
rect 447468 1300 447474 1352
rect 448422 1300 448428 1352
rect 448480 1340 448486 1352
rect 453298 1340 453304 1352
rect 448480 1312 453304 1340
rect 448480 1300 448486 1312
rect 453298 1300 453304 1312
rect 453356 1300 453362 1352
rect 458818 1300 458824 1352
rect 458876 1340 458882 1352
rect 463970 1340 463976 1352
rect 458876 1312 463976 1340
rect 458876 1300 458882 1312
rect 463970 1300 463976 1312
rect 464028 1300 464034 1352
rect 468110 1300 468116 1352
rect 468168 1340 468174 1352
rect 473078 1340 473084 1352
rect 468168 1312 473084 1340
rect 468168 1300 468174 1312
rect 473078 1300 473084 1312
rect 473136 1300 473142 1352
rect 480898 1300 480904 1352
rect 480956 1340 480962 1352
rect 486418 1340 486424 1352
rect 480956 1312 486424 1340
rect 480956 1300 480962 1312
rect 486418 1300 486424 1312
rect 486476 1300 486482 1352
rect 487798 1300 487804 1352
rect 487856 1340 487862 1352
rect 493134 1340 493140 1352
rect 487856 1312 493140 1340
rect 487856 1300 487862 1312
rect 493134 1300 493140 1312
rect 493192 1300 493198 1352
rect 497090 1300 497096 1352
rect 497148 1340 497154 1352
rect 502978 1340 502984 1352
rect 497148 1312 502984 1340
rect 497148 1300 497154 1312
rect 502978 1300 502984 1312
rect 503036 1300 503042 1352
rect 504082 1300 504088 1352
rect 504140 1340 504146 1352
rect 509694 1340 509700 1352
rect 504140 1312 509700 1340
rect 504140 1300 504146 1312
rect 509694 1300 509700 1312
rect 509752 1300 509758 1352
rect 509878 1300 509884 1352
rect 509936 1340 509942 1352
rect 515766 1340 515772 1352
rect 509936 1312 515772 1340
rect 509936 1300 509942 1312
rect 515766 1300 515772 1312
rect 515824 1300 515830 1352
rect 519170 1300 519176 1352
rect 519228 1340 519234 1352
rect 525426 1340 525432 1352
rect 519228 1312 525432 1340
rect 519228 1300 519234 1312
rect 525426 1300 525432 1312
rect 525484 1300 525490 1352
rect 526070 1300 526076 1352
rect 526128 1340 526134 1352
rect 532142 1340 532148 1352
rect 526128 1312 532148 1340
rect 526128 1300 526134 1312
rect 532142 1300 532148 1312
rect 532200 1300 532206 1352
rect 534258 1300 534264 1352
rect 534316 1340 534322 1352
rect 540422 1340 540428 1352
rect 534316 1312 540428 1340
rect 534316 1300 534322 1312
rect 540422 1300 540428 1312
rect 540480 1300 540486 1352
rect 542262 1300 542268 1352
rect 542320 1340 542326 1352
rect 549070 1340 549076 1352
rect 542320 1312 549076 1340
rect 542320 1300 542326 1312
rect 549070 1300 549076 1312
rect 549128 1300 549134 1352
rect 551646 1300 551652 1352
rect 551704 1340 551710 1352
rect 558546 1340 558552 1352
rect 551704 1312 558552 1340
rect 551704 1300 551710 1312
rect 558546 1300 558552 1312
rect 558604 1300 558610 1352
rect 560938 1300 560944 1352
rect 560996 1340 561002 1352
rect 568022 1340 568028 1352
rect 560996 1312 568028 1340
rect 560996 1300 561002 1312
rect 568022 1300 568028 1312
rect 568080 1300 568086 1352
rect 571242 1300 571248 1352
rect 571300 1340 571306 1352
rect 578602 1340 578608 1352
rect 571300 1312 578608 1340
rect 571300 1300 571306 1312
rect 578602 1300 578608 1312
rect 578660 1300 578666 1352
rect 74994 1232 75000 1284
rect 75052 1272 75058 1284
rect 77110 1272 77116 1284
rect 75052 1244 77116 1272
rect 75052 1232 75058 1244
rect 77110 1232 77116 1244
rect 77168 1232 77174 1284
rect 77386 1232 77392 1284
rect 77444 1272 77450 1284
rect 79410 1272 79416 1284
rect 77444 1244 79416 1272
rect 77444 1232 77450 1244
rect 79410 1232 79416 1244
rect 79468 1232 79474 1284
rect 82078 1232 82084 1284
rect 82136 1272 82142 1284
rect 84010 1272 84016 1284
rect 82136 1244 84016 1272
rect 82136 1232 82142 1244
rect 84010 1232 84016 1244
rect 84068 1232 84074 1284
rect 84470 1232 84476 1284
rect 84528 1272 84534 1284
rect 86402 1272 86408 1284
rect 84528 1244 86408 1272
rect 84528 1232 84534 1244
rect 86402 1232 86408 1244
rect 86460 1232 86466 1284
rect 90358 1232 90364 1284
rect 90416 1272 90422 1284
rect 92198 1272 92204 1284
rect 90416 1244 92204 1272
rect 90416 1232 90422 1244
rect 92198 1232 92204 1244
rect 92256 1232 92262 1284
rect 92750 1232 92756 1284
rect 92808 1272 92814 1284
rect 94498 1272 94504 1284
rect 92808 1244 94504 1272
rect 92808 1232 92814 1244
rect 94498 1232 94504 1244
rect 94556 1232 94562 1284
rect 98638 1232 98644 1284
rect 98696 1272 98702 1284
rect 100294 1272 100300 1284
rect 98696 1244 100300 1272
rect 98696 1232 98702 1244
rect 100294 1232 100300 1244
rect 100352 1232 100358 1284
rect 102226 1232 102232 1284
rect 102284 1272 102290 1284
rect 103790 1272 103796 1284
rect 102284 1244 103796 1272
rect 102284 1232 102290 1244
rect 103790 1232 103796 1244
rect 103848 1232 103854 1284
rect 108114 1232 108120 1284
rect 108172 1272 108178 1284
rect 109586 1272 109592 1284
rect 108172 1244 109592 1272
rect 108172 1232 108178 1244
rect 109586 1232 109592 1244
rect 109644 1232 109650 1284
rect 110506 1232 110512 1284
rect 110564 1272 110570 1284
rect 111886 1272 111892 1284
rect 110564 1244 111892 1272
rect 110564 1232 110570 1244
rect 111886 1232 111892 1244
rect 111944 1232 111950 1284
rect 115198 1232 115204 1284
rect 115256 1272 115262 1284
rect 116578 1272 116584 1284
rect 115256 1244 116584 1272
rect 115256 1232 115262 1244
rect 116578 1232 116584 1244
rect 116636 1232 116642 1284
rect 117590 1232 117596 1284
rect 117648 1272 117654 1284
rect 118878 1272 118884 1284
rect 117648 1244 118884 1272
rect 117648 1232 117654 1244
rect 118878 1232 118884 1244
rect 118936 1232 118942 1284
rect 122282 1232 122288 1284
rect 122340 1272 122346 1284
rect 123478 1272 123484 1284
rect 122340 1244 123484 1272
rect 122340 1232 122346 1244
rect 123478 1232 123484 1244
rect 123536 1232 123542 1284
rect 124674 1232 124680 1284
rect 124732 1272 124738 1284
rect 125778 1272 125784 1284
rect 124732 1244 125784 1272
rect 124732 1232 124738 1244
rect 125778 1232 125784 1244
rect 125836 1232 125842 1284
rect 128170 1232 128176 1284
rect 128228 1272 128234 1284
rect 129274 1272 129280 1284
rect 128228 1244 129280 1272
rect 128228 1232 128234 1244
rect 129274 1232 129280 1244
rect 129332 1232 129338 1284
rect 136450 1232 136456 1284
rect 136508 1272 136514 1284
rect 137370 1272 137376 1284
rect 136508 1244 137376 1272
rect 136508 1232 136514 1244
rect 137370 1232 137376 1244
rect 137428 1232 137434 1284
rect 138842 1232 138848 1284
rect 138900 1272 138906 1284
rect 139762 1272 139768 1284
rect 138900 1244 139768 1272
rect 138900 1232 138906 1244
rect 139762 1232 139768 1244
rect 139820 1232 139826 1284
rect 140038 1232 140044 1284
rect 140096 1272 140102 1284
rect 140866 1272 140872 1284
rect 140096 1244 140872 1272
rect 140096 1232 140102 1244
rect 140866 1232 140872 1244
rect 140924 1232 140930 1284
rect 281350 1232 281356 1284
rect 281408 1272 281414 1284
rect 283098 1272 283104 1284
rect 281408 1244 283104 1272
rect 281408 1232 281414 1244
rect 283098 1232 283104 1244
rect 283156 1232 283162 1284
rect 289446 1232 289452 1284
rect 289504 1272 289510 1284
rect 291378 1272 291384 1284
rect 289504 1244 291384 1272
rect 289504 1232 289510 1244
rect 291378 1232 291384 1244
rect 291436 1232 291442 1284
rect 296438 1232 296444 1284
rect 296496 1272 296502 1284
rect 298462 1272 298468 1284
rect 296496 1244 298468 1272
rect 296496 1232 296502 1244
rect 298462 1232 298468 1244
rect 298520 1232 298526 1284
rect 303338 1232 303344 1284
rect 303396 1272 303402 1284
rect 305546 1272 305552 1284
rect 303396 1244 305552 1272
rect 303396 1232 303402 1244
rect 305546 1232 305552 1244
rect 305604 1232 305610 1284
rect 312538 1232 312544 1284
rect 312596 1272 312602 1284
rect 315022 1272 315028 1284
rect 312596 1244 315028 1272
rect 312596 1232 312602 1244
rect 315022 1232 315028 1244
rect 315080 1232 315086 1284
rect 318426 1232 318432 1284
rect 318484 1272 318490 1284
rect 320910 1272 320916 1284
rect 318484 1244 320916 1272
rect 318484 1232 318490 1244
rect 320910 1232 320916 1244
rect 320968 1232 320974 1284
rect 324222 1232 324228 1284
rect 324280 1272 324286 1284
rect 326798 1272 326804 1284
rect 324280 1244 326804 1272
rect 324280 1232 324286 1244
rect 326798 1232 326804 1244
rect 326856 1232 326862 1284
rect 330018 1232 330024 1284
rect 330076 1272 330082 1284
rect 332686 1272 332692 1284
rect 330076 1244 332692 1272
rect 330076 1232 330082 1244
rect 332686 1232 332692 1244
rect 332744 1232 332750 1284
rect 334710 1232 334716 1284
rect 334768 1272 334774 1284
rect 337470 1272 337476 1284
rect 334768 1244 337476 1272
rect 334768 1232 334774 1244
rect 337470 1232 337476 1244
rect 337528 1232 337534 1284
rect 340506 1232 340512 1284
rect 340564 1272 340570 1284
rect 343358 1272 343364 1284
rect 340564 1244 343364 1272
rect 340564 1232 340570 1244
rect 343358 1232 343364 1244
rect 343416 1232 343422 1284
rect 344002 1232 344008 1284
rect 344060 1272 344066 1284
rect 346946 1272 346952 1284
rect 344060 1244 346952 1272
rect 344060 1232 344066 1244
rect 346946 1232 346952 1244
rect 347004 1232 347010 1284
rect 348602 1232 348608 1284
rect 348660 1272 348666 1284
rect 351638 1272 351644 1284
rect 348660 1244 351644 1272
rect 348660 1232 348666 1244
rect 351638 1232 351644 1244
rect 351696 1232 351702 1284
rect 352098 1232 352104 1284
rect 352156 1272 352162 1284
rect 355226 1272 355232 1284
rect 352156 1244 355232 1272
rect 352156 1232 352162 1244
rect 355226 1232 355232 1244
rect 355284 1232 355290 1284
rect 355594 1232 355600 1284
rect 355652 1272 355658 1284
rect 358722 1272 358728 1284
rect 355652 1244 358728 1272
rect 355652 1232 355658 1244
rect 358722 1232 358728 1244
rect 358780 1232 358786 1284
rect 359090 1232 359096 1284
rect 359148 1272 359154 1284
rect 362310 1272 362316 1284
rect 359148 1244 362316 1272
rect 359148 1232 359154 1244
rect 362310 1232 362316 1244
rect 362368 1232 362374 1284
rect 363690 1232 363696 1284
rect 363748 1272 363754 1284
rect 367002 1272 367008 1284
rect 363748 1244 367008 1272
rect 363748 1232 363754 1244
rect 367002 1232 367008 1244
rect 367060 1232 367066 1284
rect 372982 1232 372988 1284
rect 373040 1272 373046 1284
rect 376478 1272 376484 1284
rect 373040 1244 376484 1272
rect 373040 1232 373046 1244
rect 376478 1232 376484 1244
rect 376536 1232 376542 1284
rect 377582 1232 377588 1284
rect 377640 1272 377646 1284
rect 381170 1272 381176 1284
rect 377640 1244 381176 1272
rect 377640 1232 377646 1244
rect 381170 1232 381176 1244
rect 381228 1232 381234 1284
rect 388070 1232 388076 1284
rect 388128 1272 388134 1284
rect 391842 1272 391848 1284
rect 388128 1244 391848 1272
rect 388128 1232 388134 1244
rect 391842 1232 391848 1244
rect 391900 1232 391906 1284
rect 393866 1232 393872 1284
rect 393924 1272 393930 1284
rect 397730 1272 397736 1284
rect 393924 1244 397736 1272
rect 393924 1232 393930 1244
rect 397730 1232 397736 1244
rect 397788 1232 397794 1284
rect 398466 1232 398472 1284
rect 398524 1272 398530 1284
rect 402514 1272 402520 1284
rect 398524 1244 402520 1272
rect 398524 1232 398530 1244
rect 402514 1232 402520 1244
rect 402572 1232 402578 1284
rect 403158 1232 403164 1284
rect 403216 1272 403222 1284
rect 407206 1272 407212 1284
rect 403216 1244 407212 1272
rect 403216 1232 403222 1244
rect 407206 1232 407212 1244
rect 407264 1232 407270 1284
rect 410058 1232 410064 1284
rect 410116 1272 410122 1284
rect 414290 1272 414296 1284
rect 410116 1244 414296 1272
rect 410116 1232 410122 1244
rect 414290 1232 414296 1244
rect 414348 1232 414354 1284
rect 418246 1232 418252 1284
rect 418304 1272 418310 1284
rect 422570 1272 422576 1284
rect 418304 1244 422576 1272
rect 418304 1232 418310 1244
rect 422570 1232 422576 1244
rect 422628 1232 422634 1284
rect 424042 1232 424048 1284
rect 424100 1272 424106 1284
rect 428458 1272 428464 1284
rect 424100 1244 428464 1272
rect 424100 1232 424106 1244
rect 428458 1232 428464 1244
rect 428516 1232 428522 1284
rect 435634 1232 435640 1284
rect 435692 1272 435698 1284
rect 439958 1272 439964 1284
rect 435692 1244 439964 1272
rect 435692 1232 435698 1244
rect 439958 1232 439964 1244
rect 440016 1232 440022 1284
rect 444926 1232 444932 1284
rect 444984 1272 444990 1284
rect 449802 1272 449808 1284
rect 444984 1244 449808 1272
rect 444984 1232 444990 1244
rect 449802 1232 449808 1244
rect 449860 1232 449866 1284
rect 450722 1232 450728 1284
rect 450780 1272 450786 1284
rect 455690 1272 455696 1284
rect 450780 1244 455696 1272
rect 450780 1232 450786 1244
rect 455690 1232 455696 1244
rect 455748 1232 455754 1284
rect 456518 1232 456524 1284
rect 456576 1272 456582 1284
rect 461578 1272 461584 1284
rect 456576 1244 461584 1272
rect 456576 1232 456582 1244
rect 461578 1232 461584 1244
rect 461636 1232 461642 1284
rect 462222 1232 462228 1284
rect 462280 1272 462286 1284
rect 467466 1272 467472 1284
rect 462280 1244 467472 1272
rect 462280 1232 462286 1244
rect 467466 1232 467472 1244
rect 467524 1232 467530 1284
rect 471606 1232 471612 1284
rect 471664 1272 471670 1284
rect 476574 1272 476580 1284
rect 471664 1244 476580 1272
rect 471664 1232 471670 1244
rect 476574 1232 476580 1244
rect 476632 1232 476638 1284
rect 479702 1232 479708 1284
rect 479760 1272 479766 1284
rect 484854 1272 484860 1284
rect 479760 1244 484860 1272
rect 479760 1232 479766 1244
rect 484854 1232 484860 1244
rect 484912 1232 484918 1284
rect 488994 1232 489000 1284
rect 489052 1272 489058 1284
rect 494698 1272 494704 1284
rect 489052 1244 494704 1272
rect 489052 1232 489058 1244
rect 494698 1232 494704 1244
rect 494756 1232 494762 1284
rect 498286 1232 498292 1284
rect 498344 1272 498350 1284
rect 503806 1272 503812 1284
rect 498344 1244 503812 1272
rect 498344 1232 498350 1244
rect 503806 1232 503812 1244
rect 503864 1232 503870 1284
rect 510982 1232 510988 1284
rect 511040 1272 511046 1284
rect 517146 1272 517152 1284
rect 511040 1244 517152 1272
rect 511040 1232 511046 1244
rect 517146 1232 517152 1244
rect 517204 1232 517210 1284
rect 517974 1232 517980 1284
rect 518032 1272 518038 1284
rect 523862 1272 523868 1284
rect 518032 1244 523868 1272
rect 518032 1232 518038 1244
rect 523862 1232 523868 1244
rect 523920 1232 523926 1284
rect 527266 1232 527272 1284
rect 527324 1272 527330 1284
rect 533706 1272 533712 1284
rect 527324 1244 533712 1272
rect 527324 1232 527330 1244
rect 533706 1232 533712 1244
rect 533764 1232 533770 1284
rect 543458 1232 543464 1284
rect 543516 1272 543522 1284
rect 550266 1272 550272 1284
rect 543516 1244 550272 1272
rect 543516 1232 543522 1244
rect 550266 1232 550272 1244
rect 550324 1232 550330 1284
rect 550450 1232 550456 1284
rect 550508 1272 550514 1284
rect 557350 1272 557356 1284
rect 550508 1244 557356 1272
rect 550508 1232 550514 1244
rect 557350 1232 557356 1244
rect 557408 1232 557414 1284
rect 562042 1232 562048 1284
rect 562100 1272 562106 1284
rect 569126 1272 569132 1284
rect 562100 1244 569132 1272
rect 562100 1232 562106 1244
rect 569126 1232 569132 1244
rect 569184 1232 569190 1284
rect 570138 1232 570144 1284
rect 570196 1272 570202 1284
rect 577406 1272 577412 1284
rect 570196 1244 577412 1272
rect 570196 1232 570202 1244
rect 577406 1232 577412 1244
rect 577464 1232 577470 1284
rect 99834 1164 99840 1216
rect 99892 1204 99898 1216
rect 101490 1204 101496 1216
rect 99892 1176 101496 1204
rect 99892 1164 99898 1176
rect 101490 1164 101496 1176
rect 101548 1164 101554 1216
rect 114002 1164 114008 1216
rect 114060 1204 114066 1216
rect 115382 1204 115388 1216
rect 114060 1176 115388 1204
rect 114060 1164 114066 1176
rect 115382 1164 115388 1176
rect 115440 1164 115446 1216
rect 311526 1164 311532 1216
rect 311584 1204 311590 1216
rect 313826 1204 313832 1216
rect 311584 1176 313832 1204
rect 311584 1164 311590 1176
rect 313826 1164 313832 1176
rect 313884 1164 313890 1216
rect 319622 1164 319628 1216
rect 319680 1204 319686 1216
rect 322106 1204 322112 1216
rect 319680 1176 322112 1204
rect 319680 1164 319686 1176
rect 322106 1164 322112 1176
rect 322164 1164 322170 1216
rect 326614 1164 326620 1216
rect 326672 1204 326678 1216
rect 329190 1204 329196 1216
rect 326672 1176 329196 1204
rect 326672 1164 326678 1176
rect 329190 1164 329196 1176
rect 329248 1164 329254 1216
rect 331122 1164 331128 1216
rect 331180 1204 331186 1216
rect 333882 1204 333888 1216
rect 331180 1176 333888 1204
rect 331180 1164 331186 1176
rect 333882 1164 333888 1176
rect 333940 1164 333946 1216
rect 337010 1164 337016 1216
rect 337068 1204 337074 1216
rect 339862 1204 339868 1216
rect 337068 1176 339868 1204
rect 337068 1164 337074 1176
rect 339862 1164 339868 1176
rect 339920 1164 339926 1216
rect 341702 1164 341708 1216
rect 341760 1204 341766 1216
rect 344554 1204 344560 1216
rect 341760 1176 344560 1204
rect 341760 1164 341766 1176
rect 344554 1164 344560 1176
rect 344612 1164 344618 1216
rect 357894 1164 357900 1216
rect 357952 1204 357958 1216
rect 361114 1204 361120 1216
rect 357952 1176 361120 1204
rect 357952 1164 357958 1176
rect 361114 1164 361120 1176
rect 361172 1164 361178 1216
rect 364886 1164 364892 1216
rect 364944 1204 364950 1216
rect 368198 1204 368204 1216
rect 364944 1176 368204 1204
rect 364944 1164 364950 1176
rect 368198 1164 368204 1176
rect 368256 1164 368262 1216
rect 375282 1164 375288 1216
rect 375340 1204 375346 1216
rect 378870 1204 378876 1216
rect 375340 1176 378876 1204
rect 375340 1164 375346 1176
rect 378870 1164 378876 1176
rect 378928 1164 378934 1216
rect 381078 1164 381084 1216
rect 381136 1204 381142 1216
rect 384758 1204 384764 1216
rect 381136 1176 384764 1204
rect 381136 1164 381142 1176
rect 384758 1164 384764 1176
rect 384816 1164 384822 1216
rect 390370 1164 390376 1216
rect 390428 1204 390434 1216
rect 394234 1204 394240 1216
rect 390428 1176 394240 1204
rect 390428 1164 390434 1176
rect 394234 1164 394240 1176
rect 394292 1164 394298 1216
rect 400858 1164 400864 1216
rect 400916 1204 400922 1216
rect 404814 1204 404820 1216
rect 400916 1176 404820 1204
rect 400916 1164 400922 1176
rect 404814 1164 404820 1176
rect 404872 1164 404878 1216
rect 407758 1164 407764 1216
rect 407816 1204 407822 1216
rect 411898 1204 411904 1216
rect 407816 1176 411904 1204
rect 407816 1164 407822 1176
rect 411898 1164 411904 1176
rect 411956 1164 411962 1216
rect 413554 1164 413560 1216
rect 413612 1204 413618 1216
rect 417878 1204 417884 1216
rect 413612 1176 417884 1204
rect 413612 1164 413618 1176
rect 417878 1164 417884 1176
rect 417936 1164 417942 1216
rect 419350 1164 419356 1216
rect 419408 1204 419414 1216
rect 423398 1204 423404 1216
rect 419408 1176 423404 1204
rect 419408 1164 419414 1176
rect 423398 1164 423404 1176
rect 423456 1164 423462 1216
rect 426342 1164 426348 1216
rect 426400 1204 426406 1216
rect 430850 1204 430856 1216
rect 426400 1176 430856 1204
rect 426400 1164 426406 1176
rect 430850 1164 430856 1176
rect 430908 1164 430914 1216
rect 441430 1164 441436 1216
rect 441488 1204 441494 1216
rect 445846 1204 445852 1216
rect 441488 1176 445852 1204
rect 441488 1164 441494 1176
rect 445846 1164 445852 1176
rect 445904 1164 445910 1216
rect 446030 1164 446036 1216
rect 446088 1204 446094 1216
rect 450906 1204 450912 1216
rect 446088 1176 450912 1204
rect 446088 1164 446094 1176
rect 450906 1164 450912 1176
rect 450964 1164 450970 1216
rect 457622 1164 457628 1216
rect 457680 1204 457686 1216
rect 462406 1204 462412 1216
rect 457680 1176 462412 1204
rect 457680 1164 457686 1176
rect 462406 1164 462412 1176
rect 462464 1164 462470 1216
rect 465810 1164 465816 1216
rect 465868 1204 465874 1216
rect 470686 1204 470692 1216
rect 465868 1176 470692 1204
rect 465868 1164 465874 1176
rect 470686 1164 470692 1176
rect 470744 1164 470750 1216
rect 475102 1164 475108 1216
rect 475160 1204 475166 1216
rect 480530 1204 480536 1216
rect 475160 1176 480536 1204
rect 475160 1164 475166 1176
rect 480530 1164 480536 1176
rect 480588 1164 480594 1216
rect 482002 1164 482008 1216
rect 482060 1204 482066 1216
rect 487246 1204 487252 1216
rect 482060 1176 487252 1204
rect 482060 1164 482066 1176
rect 487246 1164 487252 1176
rect 487304 1164 487310 1216
rect 492490 1164 492496 1216
rect 492548 1204 492554 1216
rect 498194 1204 498200 1216
rect 492548 1176 498200 1204
rect 492548 1164 492554 1176
rect 498194 1164 498200 1176
rect 498252 1164 498258 1216
rect 505186 1164 505192 1216
rect 505244 1204 505250 1216
rect 511258 1204 511264 1216
rect 505244 1176 511264 1204
rect 505244 1164 505250 1176
rect 511258 1164 511264 1176
rect 511316 1164 511322 1216
rect 513282 1164 513288 1216
rect 513340 1204 513346 1216
rect 519538 1204 519544 1216
rect 513340 1176 519544 1204
rect 513340 1164 513346 1176
rect 519538 1164 519544 1176
rect 519596 1164 519602 1216
rect 522666 1164 522672 1216
rect 522724 1204 522730 1216
rect 529014 1204 529020 1216
rect 522724 1176 529020 1204
rect 522724 1164 522730 1176
rect 529014 1164 529020 1176
rect 529072 1164 529078 1216
rect 531866 1164 531872 1216
rect 531924 1204 531930 1216
rect 538398 1204 538404 1216
rect 531924 1176 538404 1204
rect 531924 1164 531930 1176
rect 538398 1164 538404 1176
rect 538456 1164 538462 1216
rect 540054 1164 540060 1216
rect 540112 1204 540118 1216
rect 546678 1204 546684 1216
rect 540112 1176 546684 1204
rect 540112 1164 540118 1176
rect 546678 1164 546684 1176
rect 546736 1164 546742 1216
rect 548150 1164 548156 1216
rect 548208 1204 548214 1216
rect 554958 1204 554964 1216
rect 548208 1176 554964 1204
rect 548208 1164 548214 1176
rect 554958 1164 554964 1176
rect 555016 1164 555022 1216
rect 558454 1164 558460 1216
rect 558512 1204 558518 1216
rect 565630 1204 565636 1216
rect 558512 1176 565636 1204
rect 558512 1164 558518 1176
rect 565630 1164 565636 1176
rect 565688 1164 565694 1216
rect 569034 1164 569040 1216
rect 569092 1204 569098 1216
rect 576302 1204 576308 1216
rect 569092 1176 576308 1204
rect 569092 1164 569098 1176
rect 576302 1164 576308 1176
rect 576360 1164 576366 1216
rect 5626 1096 5632 1148
rect 5684 1136 5690 1148
rect 8662 1136 8668 1148
rect 5684 1108 8668 1136
rect 5684 1096 5690 1108
rect 8662 1096 8668 1108
rect 8720 1096 8726 1148
rect 111610 1096 111616 1148
rect 111668 1136 111674 1148
rect 113082 1136 113088 1148
rect 111668 1108 113088 1136
rect 111668 1096 111674 1108
rect 113082 1096 113088 1108
rect 113140 1096 113146 1148
rect 123478 1096 123484 1148
rect 123536 1136 123542 1148
rect 124766 1136 124772 1148
rect 123536 1108 124772 1136
rect 123536 1096 123542 1108
rect 124766 1096 124772 1108
rect 124824 1096 124830 1148
rect 320818 1096 320824 1148
rect 320876 1136 320882 1148
rect 323302 1136 323308 1148
rect 320876 1108 323308 1136
rect 320876 1096 320882 1108
rect 323302 1096 323308 1108
rect 323360 1096 323366 1148
rect 327718 1096 327724 1148
rect 327776 1136 327782 1148
rect 330386 1136 330392 1148
rect 327776 1108 330392 1136
rect 327776 1096 327782 1108
rect 330386 1096 330392 1108
rect 330444 1096 330450 1148
rect 360102 1096 360108 1148
rect 360160 1136 360166 1148
rect 363506 1136 363512 1148
rect 360160 1108 363512 1136
rect 360160 1096 360166 1108
rect 363506 1096 363512 1108
rect 363564 1096 363570 1148
rect 382182 1096 382188 1148
rect 382240 1136 382246 1148
rect 385954 1136 385960 1148
rect 382240 1108 385960 1136
rect 382240 1096 382246 1108
rect 385954 1096 385960 1108
rect 386012 1096 386018 1148
rect 389266 1096 389272 1148
rect 389324 1136 389330 1148
rect 393038 1136 393044 1148
rect 389324 1108 393044 1136
rect 389324 1096 389330 1108
rect 393038 1096 393044 1108
rect 393096 1096 393102 1148
rect 397362 1096 397368 1148
rect 397420 1136 397426 1148
rect 401318 1136 401324 1148
rect 397420 1108 401324 1136
rect 397420 1096 397426 1108
rect 401318 1096 401324 1108
rect 401376 1096 401382 1148
rect 404262 1096 404268 1148
rect 404320 1136 404326 1148
rect 408402 1136 408408 1148
rect 404320 1108 408408 1136
rect 404320 1096 404326 1108
rect 408402 1096 408408 1108
rect 408460 1096 408466 1148
rect 408954 1096 408960 1148
rect 409012 1136 409018 1148
rect 413094 1136 413100 1148
rect 409012 1108 413100 1136
rect 409012 1096 409018 1108
rect 413094 1096 413100 1108
rect 413152 1096 413158 1148
rect 420546 1096 420552 1148
rect 420604 1136 420610 1148
rect 424962 1136 424968 1148
rect 420604 1108 424968 1136
rect 420604 1096 420610 1108
rect 424962 1096 424968 1108
rect 425020 1096 425026 1148
rect 428642 1096 428648 1148
rect 428700 1136 428706 1148
rect 433242 1136 433248 1148
rect 428700 1108 433248 1136
rect 428700 1096 428706 1108
rect 433242 1096 433248 1108
rect 433300 1096 433306 1148
rect 436738 1096 436744 1148
rect 436796 1136 436802 1148
rect 441522 1136 441528 1148
rect 436796 1108 441528 1136
rect 436796 1096 436802 1108
rect 441522 1096 441528 1108
rect 441580 1096 441586 1148
rect 454218 1096 454224 1148
rect 454276 1136 454282 1148
rect 459186 1136 459192 1148
rect 454276 1108 459192 1136
rect 454276 1096 454282 1108
rect 459186 1096 459192 1108
rect 459244 1096 459250 1148
rect 461118 1096 461124 1148
rect 461176 1136 461182 1148
rect 466270 1136 466276 1148
rect 461176 1108 466276 1136
rect 461176 1096 461182 1108
rect 466270 1096 466276 1108
rect 466328 1096 466334 1148
rect 472710 1096 472716 1148
rect 472768 1136 472774 1148
rect 478138 1136 478144 1148
rect 472768 1108 478144 1136
rect 472768 1096 472774 1108
rect 478138 1096 478144 1108
rect 478196 1096 478202 1148
rect 486694 1096 486700 1148
rect 486752 1136 486758 1148
rect 492306 1136 492312 1148
rect 486752 1108 492312 1136
rect 486752 1096 486758 1108
rect 492306 1096 492312 1108
rect 492364 1096 492370 1148
rect 493594 1096 493600 1148
rect 493652 1136 493658 1148
rect 499390 1136 499396 1148
rect 493652 1108 499396 1136
rect 493652 1096 493658 1108
rect 499390 1096 499396 1108
rect 499448 1096 499454 1148
rect 500494 1096 500500 1148
rect 500552 1136 500558 1148
rect 506474 1136 506480 1148
rect 500552 1108 506480 1136
rect 500552 1096 500558 1108
rect 506474 1096 506480 1108
rect 506532 1096 506538 1148
rect 512178 1096 512184 1148
rect 512236 1136 512242 1148
rect 517974 1136 517980 1148
rect 512236 1108 517980 1136
rect 512236 1096 512242 1108
rect 517974 1096 517980 1108
rect 518032 1096 518038 1148
rect 523770 1096 523776 1148
rect 523828 1136 523834 1148
rect 530118 1136 530124 1148
rect 523828 1108 530124 1136
rect 523828 1096 523834 1108
rect 530118 1096 530124 1108
rect 530176 1096 530182 1148
rect 530762 1096 530768 1148
rect 530820 1136 530826 1148
rect 537202 1136 537208 1148
rect 530820 1108 537208 1136
rect 530820 1096 530826 1108
rect 537202 1096 537208 1108
rect 537260 1096 537266 1148
rect 538858 1096 538864 1148
rect 538916 1136 538922 1148
rect 545482 1136 545488 1148
rect 538916 1108 545488 1136
rect 538916 1096 538922 1108
rect 545482 1096 545488 1108
rect 545540 1096 545546 1148
rect 552750 1096 552756 1148
rect 552808 1136 552814 1148
rect 559742 1136 559748 1148
rect 552808 1108 559748 1136
rect 552808 1096 552814 1108
rect 559742 1096 559748 1108
rect 559800 1096 559806 1148
rect 567838 1096 567844 1148
rect 567896 1136 567902 1148
rect 575106 1136 575112 1148
rect 567896 1108 575112 1136
rect 567896 1096 567902 1108
rect 575106 1096 575112 1108
rect 575164 1096 575170 1148
rect 378778 1028 378784 1080
rect 378836 1068 378842 1080
rect 382366 1068 382372 1080
rect 378836 1040 382372 1068
rect 378836 1028 378842 1040
rect 382366 1028 382372 1040
rect 382424 1028 382430 1080
rect 386874 1028 386880 1080
rect 386932 1068 386938 1080
rect 390646 1068 390652 1080
rect 386932 1040 390652 1068
rect 386932 1028 386938 1040
rect 390646 1028 390652 1040
rect 390704 1028 390710 1080
rect 425146 1028 425152 1080
rect 425204 1068 425210 1080
rect 429654 1068 429660 1080
rect 425204 1040 429660 1068
rect 425204 1028 425210 1040
rect 429654 1028 429660 1040
rect 429712 1028 429718 1080
rect 439130 1028 439136 1080
rect 439188 1068 439194 1080
rect 443822 1068 443828 1080
rect 439188 1040 443828 1068
rect 439188 1028 439194 1040
rect 443822 1028 443828 1040
rect 443880 1028 443886 1080
rect 447226 1028 447232 1080
rect 447284 1068 447290 1080
rect 452102 1068 452108 1080
rect 447284 1040 452108 1068
rect 447284 1028 447290 1040
rect 452102 1028 452108 1040
rect 452160 1028 452166 1080
rect 455322 1028 455328 1080
rect 455380 1068 455386 1080
rect 460106 1068 460112 1080
rect 455380 1040 460112 1068
rect 455380 1028 455386 1040
rect 460106 1028 460112 1040
rect 460164 1028 460170 1080
rect 466914 1028 466920 1080
rect 466972 1068 466978 1080
rect 472250 1068 472256 1080
rect 466972 1040 472256 1068
rect 466972 1028 466978 1040
rect 472250 1028 472256 1040
rect 472308 1028 472314 1080
rect 477402 1028 477408 1080
rect 477460 1068 477466 1080
rect 482462 1068 482468 1080
rect 477460 1040 482468 1068
rect 477460 1028 477466 1040
rect 482462 1028 482468 1040
rect 482520 1028 482526 1080
rect 485498 1028 485504 1080
rect 485556 1068 485562 1080
rect 490742 1068 490748 1080
rect 485556 1040 490748 1068
rect 485556 1028 485562 1040
rect 490742 1028 490748 1040
rect 490800 1028 490806 1080
rect 494790 1028 494796 1080
rect 494848 1068 494854 1080
rect 500586 1068 500592 1080
rect 494848 1040 500592 1068
rect 494848 1028 494854 1040
rect 500586 1028 500592 1040
rect 500644 1028 500650 1080
rect 501690 1028 501696 1080
rect 501748 1068 501754 1080
rect 507302 1068 507308 1080
rect 501748 1040 507308 1068
rect 501748 1028 501754 1040
rect 507302 1028 507308 1040
rect 507360 1028 507366 1080
rect 514478 1028 514484 1080
rect 514536 1068 514542 1080
rect 520734 1068 520740 1080
rect 514536 1040 520740 1068
rect 514536 1028 514542 1040
rect 520734 1028 520740 1040
rect 520792 1028 520798 1080
rect 521470 1028 521476 1080
rect 521528 1068 521534 1080
rect 527818 1068 527824 1080
rect 521528 1040 527824 1068
rect 521528 1028 521534 1040
rect 527818 1028 527824 1040
rect 527876 1028 527882 1080
rect 529566 1028 529572 1080
rect 529624 1068 529630 1080
rect 536098 1068 536104 1080
rect 529624 1040 536104 1068
rect 529624 1028 529630 1040
rect 536098 1028 536104 1040
rect 536156 1028 536162 1080
rect 549346 1028 549352 1080
rect 549404 1068 549410 1080
rect 556154 1068 556160 1080
rect 549404 1040 556160 1068
rect 549404 1028 549410 1040
rect 556154 1028 556160 1040
rect 556212 1028 556218 1080
rect 559650 1028 559656 1080
rect 559708 1068 559714 1080
rect 566826 1068 566832 1080
rect 559708 1040 566832 1068
rect 559708 1028 559714 1040
rect 566826 1028 566832 1040
rect 566884 1028 566890 1080
rect 374178 960 374184 1012
rect 374236 1000 374242 1012
rect 377674 1000 377680 1012
rect 374236 972 377680 1000
rect 374236 960 374242 972
rect 377674 960 377680 972
rect 377732 960 377738 1012
rect 379882 960 379888 1012
rect 379940 1000 379946 1012
rect 383562 1000 383568 1012
rect 379940 972 383568 1000
rect 379940 960 379946 972
rect 383562 960 383568 972
rect 383620 960 383626 1012
rect 414750 960 414756 1012
rect 414808 1000 414814 1012
rect 418982 1000 418988 1012
rect 414808 972 418988 1000
rect 414808 960 414814 972
rect 418982 960 418988 972
rect 419040 960 419046 1012
rect 422846 960 422852 1012
rect 422904 1000 422910 1012
rect 427262 1000 427268 1012
rect 422904 972 427268 1000
rect 422904 960 422910 972
rect 427262 960 427268 972
rect 427320 960 427326 1012
rect 432138 960 432144 1012
rect 432196 1000 432202 1012
rect 436738 1000 436744 1012
rect 432196 972 436744 1000
rect 432196 960 432202 972
rect 436738 960 436744 972
rect 436796 960 436802 1012
rect 453022 960 453028 1012
rect 453080 1000 453086 1012
rect 458082 1000 458088 1012
rect 453080 972 458088 1000
rect 453080 960 453086 972
rect 458082 960 458088 972
rect 458140 960 458146 1012
rect 464614 960 464620 1012
rect 464672 1000 464678 1012
rect 469858 1000 469864 1012
rect 464672 972 469864 1000
rect 464672 960 464678 972
rect 469858 960 469864 972
rect 469916 960 469922 1012
rect 473906 960 473912 1012
rect 473964 1000 473970 1012
rect 479334 1000 479340 1012
rect 473964 972 479340 1000
rect 473964 960 473970 972
rect 479334 960 479340 972
rect 479392 960 479398 1012
rect 484302 960 484308 1012
rect 484360 1000 484366 1012
rect 489914 1000 489920 1012
rect 484360 972 489920 1000
rect 484360 960 484366 972
rect 489914 960 489920 972
rect 489972 960 489978 1012
rect 490098 960 490104 1012
rect 490156 1000 490162 1012
rect 495526 1000 495532 1012
rect 490156 972 495532 1000
rect 490156 960 490162 972
rect 495526 960 495532 972
rect 495584 960 495590 1012
rect 495986 960 495992 1012
rect 496044 1000 496050 1012
rect 501782 1000 501788 1012
rect 496044 972 501788 1000
rect 496044 960 496050 972
rect 501782 960 501788 972
rect 501840 960 501846 1012
rect 502886 960 502892 1012
rect 502944 1000 502950 1012
rect 508866 1000 508872 1012
rect 502944 972 508872 1000
rect 502944 960 502950 972
rect 508866 960 508872 972
rect 508924 960 508930 1012
rect 520182 960 520188 1012
rect 520240 1000 520246 1012
rect 526622 1000 526628 1012
rect 520240 972 526628 1000
rect 520240 960 520246 972
rect 526622 960 526628 972
rect 526680 960 526686 1012
rect 533062 960 533068 1012
rect 533120 1000 533126 1012
rect 539594 1000 539600 1012
rect 533120 972 539600 1000
rect 533120 960 533126 972
rect 539594 960 539600 972
rect 539652 960 539658 1012
rect 8754 892 8760 944
rect 8812 932 8818 944
rect 12158 932 12164 944
rect 8812 904 12164 932
rect 8812 892 8818 904
rect 12158 892 12164 904
rect 12216 892 12222 944
rect 121086 892 121092 944
rect 121144 932 121150 944
rect 122374 932 122380 944
rect 121144 904 122380 932
rect 121144 892 121150 904
rect 122374 892 122380 904
rect 122432 892 122438 944
rect 437934 892 437940 944
rect 437992 932 437998 944
rect 442626 932 442632 944
rect 437992 904 442632 932
rect 437992 892 437998 904
rect 442626 892 442632 904
rect 442684 892 442690 944
rect 483198 892 483204 944
rect 483256 932 483262 944
rect 488810 932 488816 944
rect 483256 904 488816 932
rect 483256 892 483262 904
rect 488810 892 488816 904
rect 488868 892 488874 944
rect 491202 892 491208 944
rect 491260 932 491266 944
rect 497090 932 497096 944
rect 491260 904 497096 932
rect 491260 892 491266 904
rect 497090 892 497096 904
rect 497148 892 497154 944
rect 347498 824 347504 876
rect 347556 864 347562 876
rect 350442 864 350448 876
rect 347556 836 350448 864
rect 347556 824 347562 836
rect 350442 824 350448 836
rect 350500 824 350506 876
rect 361390 824 361396 876
rect 361448 864 361454 876
rect 364610 864 364616 876
rect 361448 836 364616 864
rect 361448 824 361454 836
rect 364610 824 364616 836
rect 364668 824 364674 876
rect 368382 824 368388 876
rect 368440 864 368446 876
rect 371694 864 371700 876
rect 368440 836 371700 864
rect 368440 824 368446 836
rect 371694 824 371700 836
rect 371752 824 371758 876
rect 371786 824 371792 876
rect 371844 864 371850 876
rect 375282 864 375288 876
rect 371844 836 375288 864
rect 371844 824 371850 836
rect 375282 824 375288 836
rect 375340 824 375346 876
rect 384574 824 384580 876
rect 384632 864 384638 876
rect 388254 864 388260 876
rect 384632 836 388260 864
rect 384632 824 384638 836
rect 388254 824 388260 836
rect 388312 824 388318 876
rect 391566 824 391572 876
rect 391624 864 391630 876
rect 395338 864 395344 876
rect 391624 836 395344 864
rect 391624 824 391630 836
rect 395338 824 395344 836
rect 395396 824 395402 876
rect 396166 824 396172 876
rect 396224 864 396230 876
rect 400122 864 400128 876
rect 396224 836 400128 864
rect 396224 824 396230 836
rect 400122 824 400128 836
rect 400180 824 400186 876
rect 406654 824 406660 876
rect 406712 864 406718 876
rect 410794 864 410800 876
rect 406712 836 410800 864
rect 406712 824 406718 836
rect 410794 824 410800 836
rect 410852 824 410858 876
rect 417050 824 417056 876
rect 417108 864 417114 876
rect 421374 864 421380 876
rect 417108 836 421380 864
rect 417108 824 417114 836
rect 421374 824 421380 836
rect 421432 824 421438 876
rect 429838 824 429844 876
rect 429896 864 429902 876
rect 434438 864 434444 876
rect 429896 836 434444 864
rect 429896 824 429902 836
rect 434438 824 434444 836
rect 434496 824 434502 876
rect 443730 824 443736 876
rect 443788 864 443794 876
rect 448238 864 448244 876
rect 443788 836 448244 864
rect 443788 824 443794 836
rect 448238 824 448244 836
rect 448296 824 448302 876
rect 451826 824 451832 876
rect 451884 864 451890 876
rect 456518 864 456524 876
rect 451884 836 456524 864
rect 451884 824 451890 836
rect 456518 824 456524 836
rect 456576 824 456582 876
rect 463418 824 463424 876
rect 463476 864 463482 876
rect 468662 864 468668 876
rect 463476 836 468668 864
rect 463476 824 463482 836
rect 468662 824 468668 836
rect 468720 824 468726 876
rect 476206 824 476212 876
rect 476264 864 476270 876
rect 481358 864 481364 876
rect 476264 836 481364 864
rect 476264 824 476270 836
rect 481358 824 481364 836
rect 481416 824 481422 876
rect 434346 756 434352 808
rect 434404 796 434410 808
rect 439130 796 439136 808
rect 434404 768 439136 796
rect 434404 756 434410 768
rect 439130 756 439136 768
rect 439188 756 439194 808
rect 52546 688 52552 740
rect 52604 728 52610 740
rect 55030 728 55036 740
rect 52604 700 55036 728
rect 52604 688 52610 700
rect 55030 688 55036 700
rect 55088 688 55094 740
rect 59630 688 59636 740
rect 59688 728 59694 740
rect 61930 728 61936 740
rect 59688 700 61936 728
rect 59688 688 59694 700
rect 61930 688 61936 700
rect 61988 688 61994 740
rect 105722 688 105728 740
rect 105780 728 105786 740
rect 107286 728 107292 740
rect 105780 700 107292 728
rect 105780 688 105786 700
rect 107286 688 107292 700
rect 107344 688 107350 740
rect 274358 688 274364 740
rect 274416 728 274422 740
rect 276014 728 276020 740
rect 274416 700 276020 728
rect 274416 688 274422 700
rect 276014 688 276020 700
rect 276072 688 276078 740
rect 333514 688 333520 740
rect 333572 728 333578 740
rect 336274 728 336280 740
rect 333572 700 336280 728
rect 333572 688 333578 700
rect 336274 688 336280 700
rect 336332 688 336338 740
rect 338206 688 338212 740
rect 338264 728 338270 740
rect 340966 728 340972 740
rect 338264 700 340972 728
rect 338264 688 338270 700
rect 340966 688 340972 700
rect 341024 688 341030 740
rect 342806 688 342812 740
rect 342864 728 342870 740
rect 345750 728 345756 740
rect 342864 700 345756 728
rect 342864 688 342870 700
rect 345750 688 345756 700
rect 345808 688 345814 740
rect 346302 688 346308 740
rect 346360 728 346366 740
rect 349246 728 349252 740
rect 346360 700 349252 728
rect 346360 688 346366 700
rect 349246 688 349252 700
rect 349304 688 349310 740
rect 350902 688 350908 740
rect 350960 728 350966 740
rect 354030 728 354036 740
rect 350960 700 354036 728
rect 350960 688 350966 700
rect 354030 688 354036 700
rect 354088 688 354094 740
rect 365990 688 365996 740
rect 366048 728 366054 740
rect 369394 728 369400 740
rect 366048 700 369400 728
rect 366048 688 366054 700
rect 369394 688 369400 700
rect 369452 688 369458 740
rect 369486 688 369492 740
rect 369544 728 369550 740
rect 372890 728 372896 740
rect 369544 700 372896 728
rect 369544 688 369550 700
rect 372890 688 372896 700
rect 372948 688 372954 740
rect 541158 688 541164 740
rect 541216 728 541222 740
rect 547874 728 547880 740
rect 541216 700 547880 728
rect 541216 688 541222 700
rect 547874 688 547880 700
rect 547932 688 547938 740
rect 557534 688 557540 740
rect 557592 728 557598 740
rect 564434 728 564440 740
rect 557592 700 564440 728
rect 557592 688 557598 700
rect 564434 688 564440 700
rect 564492 688 564498 740
rect 553946 620 553952 672
rect 554004 660 554010 672
rect 554004 632 557534 660
rect 554004 620 554010 632
rect 69106 552 69112 604
rect 69164 592 69170 604
rect 71314 592 71320 604
rect 69164 564 71320 592
rect 69164 552 69170 564
rect 71314 552 71320 564
rect 71372 552 71378 604
rect 290642 552 290648 604
rect 290700 592 290706 604
rect 292574 592 292580 604
rect 290700 564 292580 592
rect 290700 552 290706 564
rect 292574 552 292580 564
rect 292632 552 292638 604
rect 304534 552 304540 604
rect 304592 592 304598 604
rect 306742 592 306748 604
rect 304592 564 306748 592
rect 304592 552 304598 564
rect 306742 552 306748 564
rect 306800 552 306806 604
rect 556246 552 556252 604
rect 556304 552 556310 604
rect 557506 592 557534 632
rect 563146 620 563152 672
rect 563204 660 563210 672
rect 570322 660 570328 672
rect 563204 632 570328 660
rect 563204 620 563210 632
rect 570322 620 570328 632
rect 570380 620 570386 672
rect 560846 592 560852 604
rect 557506 564 560852 592
rect 560846 552 560852 564
rect 560904 552 560910 604
rect 563238 552 563244 604
rect 563296 552 563302 604
rect 556264 524 556292 552
rect 563256 524 563284 552
rect 556264 496 563284 524
rect 507486 416 507492 468
rect 507544 456 507550 468
rect 513374 456 513380 468
rect 507544 428 513380 456
rect 507544 416 507550 428
rect 513374 416 513380 428
rect 513432 416 513438 468
rect 536558 416 536564 468
rect 536616 456 536622 468
rect 542814 456 542820 468
rect 536616 428 542820 456
rect 536616 416 536622 428
rect 542814 416 542820 428
rect 542872 416 542878 468
rect 544654 416 544660 468
rect 544712 456 544718 468
rect 551094 456 551100 468
rect 544712 428 551100 456
rect 544712 416 544718 428
rect 551094 416 551100 428
rect 551152 416 551158 468
rect 566642 416 566648 468
rect 566700 456 566706 468
rect 573726 456 573732 468
rect 566700 428 573732 456
rect 566700 416 566706 428
rect 573726 416 573732 428
rect 573784 416 573790 468
rect 383378 348 383384 400
rect 383436 388 383442 400
rect 386782 388 386788 400
rect 383436 360 386788 388
rect 383436 348 383442 360
rect 386782 348 386788 360
rect 386840 348 386846 400
rect 535362 348 535368 400
rect 535420 388 535426 400
rect 542170 388 542176 400
rect 535420 360 542176 388
rect 535420 348 535426 360
rect 542170 348 542176 360
rect 542228 348 542234 400
rect 546954 348 546960 400
rect 547012 388 547018 400
rect 553946 388 553952 400
rect 547012 360 553952 388
rect 547012 348 547018 360
rect 553946 348 553952 360
rect 554004 348 554010 400
rect 537662 280 537668 332
rect 537720 320 537726 332
rect 544562 320 544568 332
rect 537720 292 544568 320
rect 537720 280 537726 292
rect 544562 280 544568 292
rect 544620 280 544626 332
rect 545850 280 545856 332
rect 545908 320 545914 332
rect 552382 320 552388 332
rect 545908 292 552388 320
rect 545908 280 545914 292
rect 552382 280 552388 292
rect 552440 280 552446 332
rect 573634 280 573640 332
rect 573692 320 573698 332
rect 581178 320 581184 332
rect 573692 292 581184 320
rect 573692 280 573698 292
rect 581178 280 581184 292
rect 581236 280 581242 332
rect 392670 212 392676 264
rect 392728 252 392734 264
rect 396166 252 396172 264
rect 392728 224 396172 252
rect 392728 212 392734 224
rect 396166 212 396172 224
rect 396224 212 396230 264
rect 412450 212 412456 264
rect 412508 252 412514 264
rect 416866 252 416872 264
rect 412508 224 416872 252
rect 412508 212 412514 224
rect 416866 212 416872 224
rect 416924 212 416930 264
rect 421742 212 421748 264
rect 421800 252 421806 264
rect 425790 252 425796 264
rect 421800 224 425796 252
rect 421800 212 421806 224
rect 425790 212 425796 224
rect 425848 212 425854 264
rect 469306 212 469312 264
rect 469364 252 469370 264
rect 474182 252 474188 264
rect 469364 224 474188 252
rect 469364 212 469370 224
rect 474182 212 474188 224
rect 474240 212 474246 264
rect 508682 212 508688 264
rect 508740 252 508746 264
rect 514938 252 514944 264
rect 508740 224 514944 252
rect 508740 212 508746 224
rect 514938 212 514944 224
rect 514996 212 515002 264
rect 528462 212 528468 264
rect 528520 252 528526 264
rect 534534 252 534540 264
rect 528520 224 534540 252
rect 528520 212 528526 224
rect 534534 212 534540 224
rect 534592 212 534598 264
rect 564250 144 564256 196
rect 564308 184 564314 196
rect 571334 184 571340 196
rect 564308 156 571340 184
rect 564308 144 564314 156
rect 571334 144 571340 156
rect 571392 144 571398 196
rect 574830 144 574836 196
rect 574888 184 574894 196
rect 581822 184 581828 196
rect 574888 156 581828 184
rect 574888 144 574894 156
rect 581822 144 581828 156
rect 581880 144 581886 196
rect 431034 76 431040 128
rect 431092 116 431098 128
rect 435174 116 435180 128
rect 431092 88 435180 116
rect 431092 76 431098 88
rect 435174 76 435180 88
rect 435232 76 435238 128
rect 460014 76 460020 128
rect 460072 116 460078 128
rect 464982 116 464988 128
rect 460072 88 464988 116
rect 460072 76 460078 88
rect 464982 76 464988 88
rect 465040 76 465046 128
rect 470410 76 470416 128
rect 470468 116 470474 128
rect 475930 116 475936 128
rect 470468 88 475936 116
rect 470468 76 470474 88
rect 475930 76 475936 88
rect 475988 76 475994 128
rect 515674 76 515680 128
rect 515732 116 515738 128
rect 521654 116 521660 128
rect 515732 88 521660 116
rect 515732 76 515738 88
rect 521654 76 521660 88
rect 521712 76 521718 128
rect 524966 76 524972 128
rect 525024 116 525030 128
rect 531498 116 531504 128
rect 525024 88 531504 116
rect 525024 76 525030 88
rect 531498 76 531504 88
rect 531556 76 531562 128
rect 555142 76 555148 128
rect 555200 116 555206 128
rect 562226 116 562232 128
rect 555200 88 562232 116
rect 555200 76 555206 88
rect 562226 76 562232 88
rect 562284 76 562290 128
rect 565446 76 565452 128
rect 565504 116 565510 128
rect 572898 116 572904 128
rect 565504 88 572904 116
rect 565504 76 565510 88
rect 572898 76 572904 88
rect 572956 76 572962 128
rect 576118 76 576124 128
rect 576176 116 576182 128
rect 583570 116 583576 128
rect 576176 88 583576 116
rect 576176 76 576182 88
rect 583570 76 583576 88
rect 583628 76 583634 128
rect 354398 8 354404 60
rect 354456 48 354462 60
rect 357342 48 357348 60
rect 354456 20 357348 48
rect 354456 8 354462 20
rect 357342 8 357348 20
rect 357400 8 357406 60
rect 401962 8 401968 60
rect 402020 48 402026 60
rect 406194 48 406200 60
rect 402020 20 406200 48
rect 402020 8 402026 20
rect 406194 8 406200 20
rect 406252 8 406258 60
rect 499206 8 499212 60
rect 499264 48 499270 60
rect 505554 48 505560 60
rect 499264 20 505560 48
rect 499264 8 499270 20
rect 505554 8 505560 20
rect 505612 8 505618 60
rect 506290 8 506296 60
rect 506348 48 506354 60
rect 512086 48 512092 60
rect 506348 20 512092 48
rect 506348 8 506354 20
rect 512086 8 512092 20
rect 512144 8 512150 60
rect 516778 8 516784 60
rect 516836 48 516842 60
rect 523218 48 523224 60
rect 516836 20 523224 48
rect 516836 8 516842 20
rect 523218 8 523224 20
rect 523276 8 523282 60
rect 572530 8 572536 60
rect 572588 48 572594 60
rect 579614 48 579620 60
rect 572588 20 579620 48
rect 572588 8 572594 20
rect 579614 8 579620 20
rect 579672 8 579678 60
<< via1 >>
rect 102048 700748 102100 700800
rect 105452 700748 105504 700800
rect 200028 700748 200080 700800
rect 202788 700748 202840 700800
rect 314476 700748 314528 700800
rect 316316 700748 316368 700800
rect 53012 700544 53064 700596
rect 56784 700544 56836 700596
rect 151084 700544 151136 700596
rect 154120 700544 154172 700596
rect 412456 700408 412508 700460
rect 413652 700408 413704 700460
rect 363512 700340 363564 700392
rect 364984 700340 365036 700392
rect 20352 700204 20404 700256
rect 24308 700204 24360 700256
rect 36728 700204 36780 700256
rect 40500 700204 40552 700256
rect 69388 700204 69440 700256
rect 72976 700204 73028 700256
rect 85764 700204 85816 700256
rect 89168 700204 89220 700256
rect 134708 700204 134760 700256
rect 137836 700204 137888 700256
rect 167368 700204 167420 700256
rect 170312 700204 170364 700256
rect 183744 700204 183796 700256
rect 186504 700204 186556 700256
rect 232780 700204 232832 700256
rect 235172 700204 235224 700256
rect 249064 700204 249116 700256
rect 251456 700204 251508 700256
rect 265440 700204 265492 700256
rect 267648 700204 267700 700256
rect 281816 700204 281868 700256
rect 283840 700204 283892 700256
rect 330760 700204 330812 700256
rect 332508 700204 332560 700256
rect 347136 700204 347188 700256
rect 348792 700204 348844 700256
rect 396172 700204 396224 700256
rect 397460 700204 397512 700256
rect 428832 700204 428884 700256
rect 429844 700204 429896 700256
rect 445208 700204 445260 700256
rect 446128 700204 446180 700256
rect 461492 700204 461544 700256
rect 462320 700204 462372 700256
rect 118424 700136 118476 700188
rect 121644 700136 121696 700188
rect 216404 700136 216456 700188
rect 218980 700136 219032 700188
rect 298008 700136 298060 700188
rect 300124 700136 300176 700188
rect 477868 700136 477920 700188
rect 478512 700136 478564 700188
rect 494244 700136 494296 700188
rect 494796 700136 494848 700188
rect 379796 699864 379848 699916
rect 381176 699864 381228 699916
rect 576768 698232 576820 698284
rect 580172 698232 580224 698284
rect 4020 698164 4072 698216
rect 8116 698164 8168 698216
rect 578332 644512 578384 644564
rect 580908 644512 580960 644564
rect 578884 257796 578936 257848
rect 580908 257796 580960 257848
rect 578516 151444 578568 151496
rect 580908 151444 580960 151496
rect 578332 44956 578384 45008
rect 579988 44956 580040 45008
rect 576860 5516 576912 5568
rect 579620 5516 579672 5568
rect 11152 3884 11204 3936
rect 14508 3884 14560 3936
rect 14740 3884 14792 3936
rect 18004 3884 18056 3936
rect 20628 3884 20680 3936
rect 23800 3884 23852 3936
rect 24216 3884 24268 3936
rect 27296 3884 27348 3936
rect 27712 3884 27764 3936
rect 30700 3884 30752 3936
rect 32404 3884 32456 3936
rect 35392 3884 35444 3936
rect 38384 3884 38436 3936
rect 41188 3884 41240 3936
rect 43076 3884 43128 3936
rect 45788 3884 45840 3936
rect 46664 3884 46716 3936
rect 49284 3884 49336 3936
rect 50160 3884 50212 3936
rect 52780 3884 52832 3936
rect 56048 3884 56100 3936
rect 58576 3884 58628 3936
rect 72608 3884 72660 3936
rect 74860 3884 74912 3936
rect 247636 3884 247688 3936
rect 248604 3884 248656 3936
rect 285908 3884 285960 3936
rect 287796 3884 287848 3936
rect 1676 3816 1728 3868
rect 5216 3816 5268 3868
rect 13544 3816 13596 3868
rect 16808 3816 16860 3868
rect 19432 3816 19484 3868
rect 22604 3816 22656 3868
rect 23020 3816 23072 3868
rect 26100 3816 26152 3868
rect 26516 3816 26568 3868
rect 29596 3816 29648 3868
rect 30104 3816 30156 3868
rect 33092 3816 33144 3868
rect 33600 3816 33652 3868
rect 36588 3816 36640 3868
rect 37188 3816 37240 3868
rect 39992 3816 40044 3868
rect 41880 3816 41932 3868
rect 44684 3816 44736 3868
rect 45468 3816 45520 3868
rect 48180 3816 48232 3868
rect 48964 3816 49016 3868
rect 51584 3816 51636 3868
rect 53748 3816 53800 3868
rect 56276 3816 56328 3868
rect 57244 3816 57296 3868
rect 59772 3816 59824 3868
rect 71504 3816 71556 3868
rect 73664 3816 73716 3868
rect 78588 3816 78640 3868
rect 80656 3816 80708 3868
rect 80888 3816 80940 3868
rect 82956 3816 83008 3868
rect 87972 3816 88024 3868
rect 89948 3816 90000 3868
rect 96252 3816 96304 3868
rect 98044 3816 98096 3868
rect 244140 3816 244192 3868
rect 245200 3816 245252 3868
rect 256928 3816 256980 3868
rect 258264 3816 258316 3868
rect 259228 3816 259280 3868
rect 260656 3816 260708 3868
rect 261620 3816 261672 3868
rect 262956 3816 263008 3868
rect 263920 3816 263972 3868
rect 265348 3816 265400 3868
rect 268520 3816 268572 3868
rect 270040 3816 270092 3868
rect 270820 3816 270872 3868
rect 272432 3816 272484 3868
rect 275512 3816 275564 3868
rect 277124 3816 277176 3868
rect 277812 3816 277864 3868
rect 279516 3816 279568 3868
rect 284804 3816 284856 3868
rect 286600 3816 286652 3868
rect 292900 3816 292952 3868
rect 294880 3816 294932 3868
rect 299892 3816 299944 3868
rect 301964 3816 302016 3868
rect 306792 3816 306844 3868
rect 309048 3816 309100 3868
rect 572 3748 624 3800
rect 4112 3748 4164 3800
rect 7656 3748 7708 3800
rect 11012 3748 11064 3800
rect 12348 3748 12400 3800
rect 15704 3748 15756 3800
rect 15936 3748 15988 3800
rect 19108 3748 19160 3800
rect 21824 3748 21876 3800
rect 24904 3748 24956 3800
rect 25320 3748 25372 3800
rect 28400 3748 28452 3800
rect 31300 3748 31352 3800
rect 34196 3748 34248 3800
rect 34796 3748 34848 3800
rect 37692 3748 37744 3800
rect 40684 3748 40736 3800
rect 43488 3748 43540 3800
rect 44272 3748 44324 3800
rect 46984 3748 47036 3800
rect 47860 3748 47912 3800
rect 50480 3748 50532 3800
rect 51356 3748 51408 3800
rect 53976 3748 54028 3800
rect 54944 3748 54996 3800
rect 57380 3748 57432 3800
rect 58440 3748 58492 3800
rect 60876 3748 60928 3800
rect 64328 3748 64380 3800
rect 66672 3748 66724 3800
rect 67088 3748 67140 3800
rect 69064 3748 69116 3800
rect 70308 3748 70360 3800
rect 72468 3748 72520 3800
rect 73804 3748 73856 3800
rect 75964 3748 76016 3800
rect 79692 3748 79744 3800
rect 81760 3748 81812 3800
rect 86868 3748 86920 3800
rect 88752 3748 88804 3800
rect 95148 3748 95200 3800
rect 96848 3748 96900 3800
rect 103336 3748 103388 3800
rect 104944 3748 104996 3800
rect 216356 3748 216408 3800
rect 216864 3748 216916 3800
rect 222152 3748 222204 3800
rect 222752 3748 222804 3800
rect 224452 3748 224504 3800
rect 225144 3748 225196 3800
rect 230248 3748 230300 3800
rect 231032 3748 231084 3800
rect 231444 3748 231496 3800
rect 232228 3748 232280 3800
rect 232548 3748 232600 3800
rect 233424 3748 233476 3800
rect 233744 3748 233796 3800
rect 234620 3748 234672 3800
rect 237240 3748 237292 3800
rect 238116 3748 238168 3800
rect 238344 3748 238396 3800
rect 239312 3748 239364 3800
rect 239540 3748 239592 3800
rect 240508 3748 240560 3800
rect 240736 3748 240788 3800
rect 241704 3748 241756 3800
rect 241840 3748 241892 3800
rect 242900 3748 242952 3800
rect 245336 3748 245388 3800
rect 246396 3748 246448 3800
rect 246532 3748 246584 3800
rect 247592 3748 247644 3800
rect 250028 3748 250080 3800
rect 251180 3748 251232 3800
rect 252328 3748 252380 3800
rect 253480 3748 253532 3800
rect 255824 3748 255876 3800
rect 257068 3748 257120 3800
rect 258124 3748 258176 3800
rect 259460 3748 259512 3800
rect 260424 3748 260476 3800
rect 261760 3748 261812 3800
rect 262724 3748 262776 3800
rect 264152 3748 264204 3800
rect 265024 3748 265076 3800
rect 266544 3748 266596 3800
rect 267416 3748 267468 3800
rect 268844 3748 268896 3800
rect 269716 3748 269768 3800
rect 271236 3748 271288 3800
rect 272016 3748 272068 3800
rect 273628 3748 273680 3800
rect 276708 3748 276760 3800
rect 278320 3748 278372 3800
rect 279008 3748 279060 3800
rect 280712 3748 280764 3800
rect 283608 3748 283660 3800
rect 285404 3748 285456 3800
rect 287104 3748 287156 3800
rect 288992 3748 289044 3800
rect 291704 3748 291756 3800
rect 293684 3748 293736 3800
rect 294096 3748 294148 3800
rect 296076 3748 296128 3800
rect 298696 3748 298748 3800
rect 300768 3748 300820 3800
rect 300996 3748 301048 3800
rect 303160 3748 303212 3800
rect 307988 3748 308040 3800
rect 310244 3748 310296 3800
rect 316084 3748 316136 3800
rect 318524 3748 318576 3800
rect 323076 3748 323128 3800
rect 325608 3748 325660 3800
rect 6460 3000 6512 3052
rect 9864 3000 9916 3052
rect 63224 3000 63276 3052
rect 65524 3000 65576 3052
rect 18236 2864 18288 2916
rect 21456 2864 21508 2916
rect 253388 2864 253440 2916
rect 254676 2864 254728 2916
rect 4068 2796 4120 2848
rect 7472 2796 7524 2848
rect 9956 2796 10008 2848
rect 13268 2796 13320 2848
rect 17040 2796 17092 2848
rect 20260 2796 20312 2848
rect 28908 2796 28960 2848
rect 31852 2796 31904 2848
rect 35992 2796 36044 2848
rect 38844 2796 38896 2848
rect 39580 2796 39632 2848
rect 42340 2796 42392 2848
rect 62028 2796 62080 2848
rect 64420 2796 64472 2848
rect 65524 2796 65576 2848
rect 67824 2796 67876 2848
rect 248880 2796 248932 2848
rect 249984 2796 250036 2848
rect 251088 2796 251140 2848
rect 252376 2796 252428 2848
rect 254584 2796 254636 2848
rect 255872 2796 255924 2848
rect 309232 2796 309284 2848
rect 311440 2796 311492 2848
rect 315028 2796 315080 2848
rect 317328 2796 317380 2848
rect 411168 2796 411220 2848
rect 415492 2796 415544 2848
rect 440148 2796 440200 2848
rect 445024 2796 445076 2848
rect 449532 2796 449584 2848
rect 454500 2796 454552 2848
rect 478512 2796 478564 2848
rect 484032 2796 484084 2848
rect 3240 1300 3292 1352
rect 6368 1300 6420 1352
rect 60832 1300 60884 1352
rect 63316 1300 63368 1352
rect 67916 1300 67968 1352
rect 70124 1300 70176 1352
rect 76196 1300 76248 1352
rect 78220 1300 78272 1352
rect 83280 1300 83332 1352
rect 85212 1300 85264 1352
rect 85672 1300 85724 1352
rect 87512 1300 87564 1352
rect 89168 1300 89220 1352
rect 91008 1300 91060 1352
rect 91560 1300 91612 1352
rect 93308 1300 93360 1352
rect 93952 1300 94004 1352
rect 95700 1300 95752 1352
rect 97448 1300 97500 1352
rect 99104 1300 99156 1352
rect 101036 1300 101088 1352
rect 102600 1300 102652 1352
rect 104532 1300 104584 1352
rect 106096 1300 106148 1352
rect 106924 1300 106976 1352
rect 108396 1300 108448 1352
rect 109316 1300 109368 1352
rect 110696 1300 110748 1352
rect 112812 1300 112864 1352
rect 114192 1300 114244 1352
rect 116400 1300 116452 1352
rect 117688 1300 117740 1352
rect 119896 1300 119948 1352
rect 121184 1300 121236 1352
rect 125876 1300 125928 1352
rect 126980 1300 127032 1352
rect 129372 1300 129424 1352
rect 130476 1300 130528 1352
rect 130568 1300 130620 1352
rect 131580 1300 131632 1352
rect 131764 1300 131816 1352
rect 132776 1300 132828 1352
rect 132960 1300 133012 1352
rect 133972 1300 134024 1352
rect 137652 1300 137704 1352
rect 138572 1300 138624 1352
rect 144736 1300 144788 1352
rect 145564 1300 145616 1352
rect 145932 1300 145984 1352
rect 146668 1300 146720 1352
rect 148324 1300 148376 1352
rect 149060 1300 149112 1352
rect 154212 1300 154264 1352
rect 154856 1300 154908 1352
rect 162492 1300 162544 1352
rect 162952 1300 163004 1352
rect 266268 1300 266320 1352
rect 267740 1300 267792 1352
rect 273168 1300 273220 1352
rect 274824 1300 274876 1352
rect 280068 1300 280120 1352
rect 281908 1300 281960 1352
rect 282552 1300 282604 1352
rect 284300 1300 284352 1352
rect 288348 1300 288400 1352
rect 290188 1300 290240 1352
rect 295248 1300 295300 1352
rect 297272 1300 297324 1352
rect 297548 1300 297600 1352
rect 299664 1300 299716 1352
rect 302148 1300 302200 1352
rect 304356 1300 304408 1352
rect 305736 1300 305788 1352
rect 307944 1300 307996 1352
rect 310336 1300 310388 1352
rect 312636 1300 312688 1352
rect 313832 1300 313884 1352
rect 316224 1300 316276 1352
rect 317236 1300 317288 1352
rect 319720 1300 319772 1352
rect 321928 1300 321980 1352
rect 324412 1300 324464 1352
rect 325424 1300 325476 1352
rect 328000 1300 328052 1352
rect 328920 1300 328972 1352
rect 331588 1300 331640 1352
rect 332416 1300 332468 1352
rect 335084 1300 335136 1352
rect 335912 1300 335964 1352
rect 338672 1300 338724 1352
rect 339316 1300 339368 1352
rect 342168 1300 342220 1352
rect 345112 1300 345164 1352
rect 348056 1300 348108 1352
rect 349804 1300 349856 1352
rect 352840 1300 352892 1352
rect 353208 1300 353260 1352
rect 356336 1300 356388 1352
rect 356704 1300 356756 1352
rect 359924 1300 359976 1352
rect 362592 1300 362644 1352
rect 365812 1300 365864 1352
rect 367192 1300 367244 1352
rect 370596 1300 370648 1352
rect 370688 1300 370740 1352
rect 374092 1300 374144 1352
rect 376392 1300 376444 1352
rect 379980 1300 380032 1352
rect 385776 1300 385828 1352
rect 389456 1300 389508 1352
rect 395068 1300 395120 1352
rect 398932 1300 398984 1352
rect 399668 1300 399720 1352
rect 403624 1300 403676 1352
rect 405464 1300 405516 1352
rect 409604 1300 409656 1352
rect 415952 1300 416004 1352
rect 420184 1300 420236 1352
rect 427544 1300 427596 1352
rect 431868 1300 431920 1352
rect 433248 1300 433300 1352
rect 437848 1300 437900 1352
rect 442632 1300 442684 1352
rect 447416 1300 447468 1352
rect 448428 1300 448480 1352
rect 453304 1300 453356 1352
rect 458824 1300 458876 1352
rect 463976 1300 464028 1352
rect 468116 1300 468168 1352
rect 473084 1300 473136 1352
rect 480904 1300 480956 1352
rect 486424 1300 486476 1352
rect 487804 1300 487856 1352
rect 493140 1300 493192 1352
rect 497096 1300 497148 1352
rect 502984 1300 503036 1352
rect 504088 1300 504140 1352
rect 509700 1300 509752 1352
rect 509884 1300 509936 1352
rect 515772 1300 515824 1352
rect 519176 1300 519228 1352
rect 525432 1300 525484 1352
rect 526076 1300 526128 1352
rect 532148 1300 532200 1352
rect 534264 1300 534316 1352
rect 540428 1300 540480 1352
rect 542268 1300 542320 1352
rect 549076 1300 549128 1352
rect 551652 1300 551704 1352
rect 558552 1300 558604 1352
rect 560944 1300 560996 1352
rect 568028 1300 568080 1352
rect 571248 1300 571300 1352
rect 578608 1300 578660 1352
rect 75000 1232 75052 1284
rect 77116 1232 77168 1284
rect 77392 1232 77444 1284
rect 79416 1232 79468 1284
rect 82084 1232 82136 1284
rect 84016 1232 84068 1284
rect 84476 1232 84528 1284
rect 86408 1232 86460 1284
rect 90364 1232 90416 1284
rect 92204 1232 92256 1284
rect 92756 1232 92808 1284
rect 94504 1232 94556 1284
rect 98644 1232 98696 1284
rect 100300 1232 100352 1284
rect 102232 1232 102284 1284
rect 103796 1232 103848 1284
rect 108120 1232 108172 1284
rect 109592 1232 109644 1284
rect 110512 1232 110564 1284
rect 111892 1232 111944 1284
rect 115204 1232 115256 1284
rect 116584 1232 116636 1284
rect 117596 1232 117648 1284
rect 118884 1232 118936 1284
rect 122288 1232 122340 1284
rect 123484 1232 123536 1284
rect 124680 1232 124732 1284
rect 125784 1232 125836 1284
rect 128176 1232 128228 1284
rect 129280 1232 129332 1284
rect 136456 1232 136508 1284
rect 137376 1232 137428 1284
rect 138848 1232 138900 1284
rect 139768 1232 139820 1284
rect 140044 1232 140096 1284
rect 140872 1232 140924 1284
rect 281356 1232 281408 1284
rect 283104 1232 283156 1284
rect 289452 1232 289504 1284
rect 291384 1232 291436 1284
rect 296444 1232 296496 1284
rect 298468 1232 298520 1284
rect 303344 1232 303396 1284
rect 305552 1232 305604 1284
rect 312544 1232 312596 1284
rect 315028 1232 315080 1284
rect 318432 1232 318484 1284
rect 320916 1232 320968 1284
rect 324228 1232 324280 1284
rect 326804 1232 326856 1284
rect 330024 1232 330076 1284
rect 332692 1232 332744 1284
rect 334716 1232 334768 1284
rect 337476 1232 337528 1284
rect 340512 1232 340564 1284
rect 343364 1232 343416 1284
rect 344008 1232 344060 1284
rect 346952 1232 347004 1284
rect 348608 1232 348660 1284
rect 351644 1232 351696 1284
rect 352104 1232 352156 1284
rect 355232 1232 355284 1284
rect 355600 1232 355652 1284
rect 358728 1232 358780 1284
rect 359096 1232 359148 1284
rect 362316 1232 362368 1284
rect 363696 1232 363748 1284
rect 367008 1232 367060 1284
rect 372988 1232 373040 1284
rect 376484 1232 376536 1284
rect 377588 1232 377640 1284
rect 381176 1232 381228 1284
rect 388076 1232 388128 1284
rect 391848 1232 391900 1284
rect 393872 1232 393924 1284
rect 397736 1232 397788 1284
rect 398472 1232 398524 1284
rect 402520 1232 402572 1284
rect 403164 1232 403216 1284
rect 407212 1232 407264 1284
rect 410064 1232 410116 1284
rect 414296 1232 414348 1284
rect 418252 1232 418304 1284
rect 422576 1232 422628 1284
rect 424048 1232 424100 1284
rect 428464 1232 428516 1284
rect 435640 1232 435692 1284
rect 439964 1232 440016 1284
rect 444932 1232 444984 1284
rect 449808 1232 449860 1284
rect 450728 1232 450780 1284
rect 455696 1232 455748 1284
rect 456524 1232 456576 1284
rect 461584 1232 461636 1284
rect 462228 1232 462280 1284
rect 467472 1232 467524 1284
rect 471612 1232 471664 1284
rect 476580 1232 476632 1284
rect 479708 1232 479760 1284
rect 484860 1232 484912 1284
rect 489000 1232 489052 1284
rect 494704 1232 494756 1284
rect 498292 1232 498344 1284
rect 503812 1232 503864 1284
rect 510988 1232 511040 1284
rect 517152 1232 517204 1284
rect 517980 1232 518032 1284
rect 523868 1232 523920 1284
rect 527272 1232 527324 1284
rect 533712 1232 533764 1284
rect 543464 1232 543516 1284
rect 550272 1232 550324 1284
rect 550456 1232 550508 1284
rect 557356 1232 557408 1284
rect 562048 1232 562100 1284
rect 569132 1232 569184 1284
rect 570144 1232 570196 1284
rect 577412 1232 577464 1284
rect 99840 1164 99892 1216
rect 101496 1164 101548 1216
rect 114008 1164 114060 1216
rect 115388 1164 115440 1216
rect 311532 1164 311584 1216
rect 313832 1164 313884 1216
rect 319628 1164 319680 1216
rect 322112 1164 322164 1216
rect 326620 1164 326672 1216
rect 329196 1164 329248 1216
rect 331128 1164 331180 1216
rect 333888 1164 333940 1216
rect 337016 1164 337068 1216
rect 339868 1164 339920 1216
rect 341708 1164 341760 1216
rect 344560 1164 344612 1216
rect 357900 1164 357952 1216
rect 361120 1164 361172 1216
rect 364892 1164 364944 1216
rect 368204 1164 368256 1216
rect 375288 1164 375340 1216
rect 378876 1164 378928 1216
rect 381084 1164 381136 1216
rect 384764 1164 384816 1216
rect 390376 1164 390428 1216
rect 394240 1164 394292 1216
rect 400864 1164 400916 1216
rect 404820 1164 404872 1216
rect 407764 1164 407816 1216
rect 411904 1164 411956 1216
rect 413560 1164 413612 1216
rect 417884 1164 417936 1216
rect 419356 1164 419408 1216
rect 423404 1164 423456 1216
rect 426348 1164 426400 1216
rect 430856 1164 430908 1216
rect 441436 1164 441488 1216
rect 445852 1164 445904 1216
rect 446036 1164 446088 1216
rect 450912 1164 450964 1216
rect 457628 1164 457680 1216
rect 462412 1164 462464 1216
rect 465816 1164 465868 1216
rect 470692 1164 470744 1216
rect 475108 1164 475160 1216
rect 480536 1164 480588 1216
rect 482008 1164 482060 1216
rect 487252 1164 487304 1216
rect 492496 1164 492548 1216
rect 498200 1164 498252 1216
rect 505192 1164 505244 1216
rect 511264 1164 511316 1216
rect 513288 1164 513340 1216
rect 519544 1164 519596 1216
rect 522672 1164 522724 1216
rect 529020 1164 529072 1216
rect 531872 1164 531924 1216
rect 538404 1164 538456 1216
rect 540060 1164 540112 1216
rect 546684 1164 546736 1216
rect 548156 1164 548208 1216
rect 554964 1164 555016 1216
rect 558460 1164 558512 1216
rect 565636 1164 565688 1216
rect 569040 1164 569092 1216
rect 576308 1164 576360 1216
rect 5632 1096 5684 1148
rect 8668 1096 8720 1148
rect 111616 1096 111668 1148
rect 113088 1096 113140 1148
rect 123484 1096 123536 1148
rect 124772 1096 124824 1148
rect 320824 1096 320876 1148
rect 323308 1096 323360 1148
rect 327724 1096 327776 1148
rect 330392 1096 330444 1148
rect 360108 1096 360160 1148
rect 363512 1096 363564 1148
rect 382188 1096 382240 1148
rect 385960 1096 386012 1148
rect 389272 1096 389324 1148
rect 393044 1096 393096 1148
rect 397368 1096 397420 1148
rect 401324 1096 401376 1148
rect 404268 1096 404320 1148
rect 408408 1096 408460 1148
rect 408960 1096 409012 1148
rect 413100 1096 413152 1148
rect 420552 1096 420604 1148
rect 424968 1096 425020 1148
rect 428648 1096 428700 1148
rect 433248 1096 433300 1148
rect 436744 1096 436796 1148
rect 441528 1096 441580 1148
rect 454224 1096 454276 1148
rect 459192 1096 459244 1148
rect 461124 1096 461176 1148
rect 466276 1096 466328 1148
rect 472716 1096 472768 1148
rect 478144 1096 478196 1148
rect 486700 1096 486752 1148
rect 492312 1096 492364 1148
rect 493600 1096 493652 1148
rect 499396 1096 499448 1148
rect 500500 1096 500552 1148
rect 506480 1096 506532 1148
rect 512184 1096 512236 1148
rect 517980 1096 518032 1148
rect 523776 1096 523828 1148
rect 530124 1096 530176 1148
rect 530768 1096 530820 1148
rect 537208 1096 537260 1148
rect 538864 1096 538916 1148
rect 545488 1096 545540 1148
rect 552756 1096 552808 1148
rect 559748 1096 559800 1148
rect 567844 1096 567896 1148
rect 575112 1096 575164 1148
rect 378784 1028 378836 1080
rect 382372 1028 382424 1080
rect 386880 1028 386932 1080
rect 390652 1028 390704 1080
rect 425152 1028 425204 1080
rect 429660 1028 429712 1080
rect 439136 1028 439188 1080
rect 443828 1028 443880 1080
rect 447232 1028 447284 1080
rect 452108 1028 452160 1080
rect 455328 1028 455380 1080
rect 460112 1028 460164 1080
rect 466920 1028 466972 1080
rect 472256 1028 472308 1080
rect 477408 1028 477460 1080
rect 482468 1028 482520 1080
rect 485504 1028 485556 1080
rect 490748 1028 490800 1080
rect 494796 1028 494848 1080
rect 500592 1028 500644 1080
rect 501696 1028 501748 1080
rect 507308 1028 507360 1080
rect 514484 1028 514536 1080
rect 520740 1028 520792 1080
rect 521476 1028 521528 1080
rect 527824 1028 527876 1080
rect 529572 1028 529624 1080
rect 536104 1028 536156 1080
rect 549352 1028 549404 1080
rect 556160 1028 556212 1080
rect 559656 1028 559708 1080
rect 566832 1028 566884 1080
rect 374184 960 374236 1012
rect 377680 960 377732 1012
rect 379888 960 379940 1012
rect 383568 960 383620 1012
rect 414756 960 414808 1012
rect 418988 960 419040 1012
rect 422852 960 422904 1012
rect 427268 960 427320 1012
rect 432144 960 432196 1012
rect 436744 960 436796 1012
rect 453028 960 453080 1012
rect 458088 960 458140 1012
rect 464620 960 464672 1012
rect 469864 960 469916 1012
rect 473912 960 473964 1012
rect 479340 960 479392 1012
rect 484308 960 484360 1012
rect 489920 960 489972 1012
rect 490104 960 490156 1012
rect 495532 960 495584 1012
rect 495992 960 496044 1012
rect 501788 960 501840 1012
rect 502892 960 502944 1012
rect 508872 960 508924 1012
rect 520188 960 520240 1012
rect 526628 960 526680 1012
rect 533068 960 533120 1012
rect 539600 960 539652 1012
rect 8760 892 8812 944
rect 12164 892 12216 944
rect 121092 892 121144 944
rect 122380 892 122432 944
rect 437940 892 437992 944
rect 442632 892 442684 944
rect 483204 892 483256 944
rect 488816 892 488868 944
rect 491208 892 491260 944
rect 497096 892 497148 944
rect 347504 824 347556 876
rect 350448 824 350500 876
rect 361396 824 361448 876
rect 364616 824 364668 876
rect 368388 824 368440 876
rect 371700 824 371752 876
rect 371792 824 371844 876
rect 375288 824 375340 876
rect 384580 824 384632 876
rect 388260 824 388312 876
rect 391572 824 391624 876
rect 395344 824 395396 876
rect 396172 824 396224 876
rect 400128 824 400180 876
rect 406660 824 406712 876
rect 410800 824 410852 876
rect 417056 824 417108 876
rect 421380 824 421432 876
rect 429844 824 429896 876
rect 434444 824 434496 876
rect 443736 824 443788 876
rect 448244 824 448296 876
rect 451832 824 451884 876
rect 456524 824 456576 876
rect 463424 824 463476 876
rect 468668 824 468720 876
rect 476212 824 476264 876
rect 481364 824 481416 876
rect 434352 756 434404 808
rect 439136 756 439188 808
rect 52552 688 52604 740
rect 55036 688 55088 740
rect 59636 688 59688 740
rect 61936 688 61988 740
rect 105728 688 105780 740
rect 107292 688 107344 740
rect 274364 688 274416 740
rect 276020 688 276072 740
rect 333520 688 333572 740
rect 336280 688 336332 740
rect 338212 688 338264 740
rect 340972 688 341024 740
rect 342812 688 342864 740
rect 345756 688 345808 740
rect 346308 688 346360 740
rect 349252 688 349304 740
rect 350908 688 350960 740
rect 354036 688 354088 740
rect 365996 688 366048 740
rect 369400 688 369452 740
rect 369492 688 369544 740
rect 372896 688 372948 740
rect 541164 688 541216 740
rect 547880 688 547932 740
rect 557540 688 557592 740
rect 564440 688 564492 740
rect 553952 620 554004 672
rect 69112 552 69164 604
rect 71320 552 71372 604
rect 290648 552 290700 604
rect 292580 552 292632 604
rect 304540 552 304592 604
rect 306748 552 306800 604
rect 556252 552 556304 604
rect 563152 620 563204 672
rect 570328 620 570380 672
rect 560852 552 560904 604
rect 563244 552 563296 604
rect 507492 416 507544 468
rect 513380 416 513432 468
rect 536564 416 536616 468
rect 542820 416 542872 468
rect 544660 416 544712 468
rect 551100 416 551152 468
rect 566648 416 566700 468
rect 573732 416 573784 468
rect 383384 348 383436 400
rect 386788 348 386840 400
rect 535368 348 535420 400
rect 542176 348 542228 400
rect 546960 348 547012 400
rect 553952 348 554004 400
rect 537668 280 537720 332
rect 544568 280 544620 332
rect 545856 280 545908 332
rect 552388 280 552440 332
rect 573640 280 573692 332
rect 581184 280 581236 332
rect 392676 212 392728 264
rect 396172 212 396224 264
rect 412456 212 412508 264
rect 416872 212 416924 264
rect 421748 212 421800 264
rect 425796 212 425848 264
rect 469312 212 469364 264
rect 474188 212 474240 264
rect 508688 212 508740 264
rect 514944 212 514996 264
rect 528468 212 528520 264
rect 534540 212 534592 264
rect 564256 144 564308 196
rect 571340 144 571392 196
rect 574836 144 574888 196
rect 581828 144 581880 196
rect 431040 76 431092 128
rect 435180 76 435232 128
rect 460020 76 460072 128
rect 464988 76 465040 128
rect 470416 76 470468 128
rect 475936 76 475988 128
rect 515680 76 515732 128
rect 521660 76 521712 128
rect 524972 76 525024 128
rect 531504 76 531556 128
rect 555148 76 555200 128
rect 562232 76 562284 128
rect 565452 76 565504 128
rect 572904 76 572956 128
rect 576124 76 576176 128
rect 583576 76 583628 128
rect 354404 8 354456 60
rect 357348 8 357400 60
rect 401968 8 402020 60
rect 406200 8 406252 60
rect 499212 8 499264 60
rect 505560 8 505612 60
rect 506296 8 506348 60
rect 512092 8 512144 60
rect 516784 8 516836 60
rect 523224 8 523276 60
rect 572536 8 572588 60
rect 579620 8 579672 60
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510632 703582 510844 703610
rect 8128 698222 8156 703520
rect 24320 700262 24348 703520
rect 40512 700262 40540 703520
rect 56796 700602 56824 703520
rect 53012 700596 53064 700602
rect 53012 700538 53064 700544
rect 56784 700596 56836 700602
rect 56784 700538 56836 700544
rect 20352 700256 20404 700262
rect 20352 700198 20404 700204
rect 24308 700256 24360 700262
rect 24308 700198 24360 700204
rect 36728 700256 36780 700262
rect 36728 700198 36780 700204
rect 40500 700256 40552 700262
rect 40500 700198 40552 700204
rect 4020 698216 4072 698222
rect 4020 698158 4072 698164
rect 8116 698216 8168 698222
rect 20364 698170 20392 700198
rect 36740 698170 36768 700198
rect 53024 698170 53052 700538
rect 72988 700262 73016 703520
rect 89180 700262 89208 703520
rect 105464 700806 105492 703520
rect 102048 700800 102100 700806
rect 102048 700742 102100 700748
rect 105452 700800 105504 700806
rect 105452 700742 105504 700748
rect 69388 700256 69440 700262
rect 69388 700198 69440 700204
rect 72976 700256 73028 700262
rect 72976 700198 73028 700204
rect 85764 700256 85816 700262
rect 85764 700198 85816 700204
rect 89168 700256 89220 700262
rect 89168 700198 89220 700204
rect 69400 698170 69428 700198
rect 85776 698170 85804 700198
rect 102060 698170 102088 700742
rect 121656 700194 121684 703520
rect 137848 700262 137876 703520
rect 154132 700602 154160 703520
rect 151084 700596 151136 700602
rect 151084 700538 151136 700544
rect 154120 700596 154172 700602
rect 154120 700538 154172 700544
rect 134708 700256 134760 700262
rect 134708 700198 134760 700204
rect 137836 700256 137888 700262
rect 137836 700198 137888 700204
rect 118424 700188 118476 700194
rect 118424 700130 118476 700136
rect 121644 700188 121696 700194
rect 121644 700130 121696 700136
rect 118436 698170 118464 700130
rect 134720 698170 134748 700198
rect 151096 698170 151124 700538
rect 170324 700262 170352 703520
rect 186516 700262 186544 703520
rect 202800 700806 202828 703520
rect 200028 700800 200080 700806
rect 200028 700742 200080 700748
rect 202788 700800 202840 700806
rect 202788 700742 202840 700748
rect 167368 700256 167420 700262
rect 167368 700198 167420 700204
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 183744 700256 183796 700262
rect 183744 700198 183796 700204
rect 186504 700256 186556 700262
rect 186504 700198 186556 700204
rect 167380 698170 167408 700198
rect 183756 698170 183784 700198
rect 8116 698158 8168 698164
rect 3514 697976 3570 697985
rect 4032 697959 4060 698158
rect 20316 698142 20392 698170
rect 36692 698142 36768 698170
rect 52976 698142 53052 698170
rect 69352 698142 69428 698170
rect 85728 698142 85804 698170
rect 102012 698142 102088 698170
rect 118388 698142 118464 698170
rect 134672 698142 134748 698170
rect 151048 698142 151124 698170
rect 167332 698142 167408 698170
rect 183708 698142 183784 698170
rect 200040 698170 200068 700742
rect 218992 700194 219020 703520
rect 235184 700262 235212 703520
rect 251468 700262 251496 703520
rect 267660 700262 267688 703520
rect 283852 700262 283880 703520
rect 232780 700256 232832 700262
rect 232780 700198 232832 700204
rect 235172 700256 235224 700262
rect 235172 700198 235224 700204
rect 249064 700256 249116 700262
rect 249064 700198 249116 700204
rect 251456 700256 251508 700262
rect 251456 700198 251508 700204
rect 265440 700256 265492 700262
rect 265440 700198 265492 700204
rect 267648 700256 267700 700262
rect 267648 700198 267700 700204
rect 281816 700256 281868 700262
rect 281816 700198 281868 700204
rect 283840 700256 283892 700262
rect 283840 700198 283892 700204
rect 216404 700188 216456 700194
rect 216404 700130 216456 700136
rect 218980 700188 219032 700194
rect 218980 700130 219032 700136
rect 216416 698170 216444 700130
rect 232792 698170 232820 700198
rect 249076 698170 249104 700198
rect 265452 698170 265480 700198
rect 281828 698170 281856 700198
rect 300136 700194 300164 703520
rect 316328 700806 316356 703520
rect 314476 700800 314528 700806
rect 314476 700742 314528 700748
rect 316316 700800 316368 700806
rect 316316 700742 316368 700748
rect 298008 700188 298060 700194
rect 298008 700130 298060 700136
rect 300124 700188 300176 700194
rect 300124 700130 300176 700136
rect 200040 698142 200112 698170
rect 20316 697959 20344 698142
rect 36692 697959 36720 698142
rect 52976 697959 53004 698142
rect 69352 697959 69380 698142
rect 85728 697959 85756 698142
rect 102012 697959 102040 698142
rect 118388 697959 118416 698142
rect 134672 697959 134700 698142
rect 151048 697959 151076 698142
rect 167332 697959 167360 698142
rect 183708 697959 183736 698142
rect 200084 697959 200112 698142
rect 216368 698142 216444 698170
rect 232744 698142 232820 698170
rect 249028 698142 249104 698170
rect 265404 698142 265480 698170
rect 281780 698142 281856 698170
rect 298020 698170 298048 700130
rect 314488 698170 314516 700742
rect 332520 700262 332548 703520
rect 348804 700262 348832 703520
rect 364996 700398 365024 703520
rect 363512 700392 363564 700398
rect 363512 700334 363564 700340
rect 364984 700392 365036 700398
rect 364984 700334 365036 700340
rect 330760 700256 330812 700262
rect 330760 700198 330812 700204
rect 332508 700256 332560 700262
rect 332508 700198 332560 700204
rect 347136 700256 347188 700262
rect 347136 700198 347188 700204
rect 348792 700256 348844 700262
rect 348792 700198 348844 700204
rect 330772 698170 330800 700198
rect 347148 698170 347176 700198
rect 363524 698170 363552 700334
rect 381188 699922 381216 703520
rect 397472 700262 397500 703520
rect 413664 700466 413692 703520
rect 412456 700460 412508 700466
rect 412456 700402 412508 700408
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 396172 700256 396224 700262
rect 396172 700198 396224 700204
rect 397460 700256 397512 700262
rect 397460 700198 397512 700204
rect 379796 699916 379848 699922
rect 379796 699858 379848 699864
rect 381176 699916 381228 699922
rect 381176 699858 381228 699864
rect 379808 698170 379836 699858
rect 396184 698170 396212 700198
rect 412468 698170 412496 700402
rect 429856 700262 429884 703520
rect 446140 700262 446168 703520
rect 462332 700262 462360 703520
rect 428832 700256 428884 700262
rect 428832 700198 428884 700204
rect 429844 700256 429896 700262
rect 429844 700198 429896 700204
rect 445208 700256 445260 700262
rect 445208 700198 445260 700204
rect 446128 700256 446180 700262
rect 446128 700198 446180 700204
rect 461492 700256 461544 700262
rect 461492 700198 461544 700204
rect 462320 700256 462372 700262
rect 462320 700198 462372 700204
rect 428844 698170 428872 700198
rect 445220 698170 445248 700198
rect 461504 698170 461532 700198
rect 478524 700194 478552 703520
rect 494808 700194 494836 703520
rect 477868 700188 477920 700194
rect 477868 700130 477920 700136
rect 478512 700188 478564 700194
rect 478512 700130 478564 700136
rect 494244 700188 494296 700194
rect 494244 700130 494296 700136
rect 494796 700188 494848 700194
rect 494796 700130 494848 700136
rect 477880 698170 477908 700130
rect 494256 698170 494284 700130
rect 510632 699802 510660 703582
rect 510816 703474 510844 703582
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 511000 703474 511028 703520
rect 510816 703446 511028 703474
rect 527192 699802 527220 703520
rect 543476 702434 543504 703520
rect 559668 702434 559696 703520
rect 510540 699774 510660 699802
rect 526916 699774 527220 699802
rect 543200 702406 543504 702434
rect 559576 702406 559696 702434
rect 510540 698170 510568 699774
rect 526916 698170 526944 699774
rect 543200 698170 543228 702406
rect 559576 698170 559604 702406
rect 298020 698142 298092 698170
rect 216368 697959 216396 698142
rect 232744 697959 232772 698142
rect 249028 697959 249056 698142
rect 265404 697959 265432 698142
rect 281780 697959 281808 698142
rect 298064 697959 298092 698142
rect 314440 698142 314516 698170
rect 330724 698142 330800 698170
rect 347100 698142 347176 698170
rect 363476 698142 363552 698170
rect 379760 698142 379836 698170
rect 396136 698142 396212 698170
rect 412420 698142 412496 698170
rect 428796 698142 428872 698170
rect 445172 698142 445248 698170
rect 461456 698142 461532 698170
rect 477832 698142 477908 698170
rect 494208 698142 494284 698170
rect 510492 698142 510568 698170
rect 526868 698142 526944 698170
rect 543152 698142 543228 698170
rect 559528 698142 559604 698170
rect 575860 698170 575888 703520
rect 576768 698284 576820 698290
rect 576768 698226 576820 698232
rect 580172 698284 580224 698290
rect 580172 698226 580224 698232
rect 576780 698193 576808 698226
rect 576766 698184 576822 698193
rect 575860 698142 575932 698170
rect 314440 697959 314468 698142
rect 330724 697959 330752 698142
rect 347100 697959 347128 698142
rect 363476 697959 363504 698142
rect 379760 697959 379788 698142
rect 396136 697959 396164 698142
rect 412420 697959 412448 698142
rect 428796 697959 428824 698142
rect 445172 697959 445200 698142
rect 461456 697959 461484 698142
rect 477832 697959 477860 698142
rect 494208 697959 494236 698142
rect 510492 697959 510520 698142
rect 526868 697959 526896 698142
rect 543152 697959 543180 698142
rect 559528 697959 559556 698142
rect 575904 697959 575932 698142
rect 576766 698119 576822 698128
rect 3514 697911 3570 697920
rect 3528 697377 3556 697911
rect 3514 697368 3570 697377
rect 3514 697303 3570 697312
rect 580184 697241 580212 698226
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 579526 684720 579582 684729
rect 579582 684678 579660 684706
rect 579526 684655 579582 684664
rect 579632 683913 579660 684678
rect 579618 683904 579674 683913
rect 579618 683839 579674 683848
rect 578330 644600 578386 644609
rect 578330 644535 578332 644544
rect 578384 644535 578386 644544
rect 580908 644564 580960 644570
rect 578332 644506 578384 644512
rect 580908 644506 580960 644512
rect 580920 644065 580948 644506
rect 580906 644056 580962 644065
rect 580906 643991 580962 644000
rect 3422 436656 3478 436665
rect 3422 436591 3478 436600
rect 3436 436051 3464 436591
rect 3422 436042 3478 436051
rect 3422 435977 3478 435986
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 422997 3464 423535
rect 3422 422988 3478 422997
rect 3422 422923 3478 422932
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3436 409943 3464 410479
rect 3422 409934 3478 409943
rect 3422 409869 3478 409878
rect 3422 397488 3478 397497
rect 3422 397423 3478 397432
rect 3436 396889 3464 397423
rect 3422 396880 3478 396889
rect 3422 396815 3478 396824
rect 3422 384432 3478 384441
rect 3422 384367 3478 384376
rect 3436 383713 3464 384367
rect 3422 383704 3478 383713
rect 3422 383639 3478 383648
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 370659 3464 371311
rect 3422 370650 3478 370659
rect 3422 370585 3478 370594
rect 3422 358456 3478 358465
rect 3422 358391 3478 358400
rect 3436 357605 3464 358391
rect 3422 357596 3478 357605
rect 3422 357531 3478 357540
rect 579526 351928 579582 351937
rect 579526 351863 579582 351872
rect 579540 351121 579568 351863
rect 579526 351112 579582 351121
rect 579526 351047 579582 351056
rect 3422 345400 3478 345409
rect 3422 345335 3478 345344
rect 3436 344429 3464 345335
rect 3422 344420 3478 344429
rect 3422 344355 3478 344364
rect 579618 338600 579674 338609
rect 579618 338535 579674 338544
rect 579526 337920 579582 337929
rect 579632 337906 579660 338535
rect 579582 337878 579660 337906
rect 579526 337855 579582 337864
rect 3422 332344 3478 332353
rect 3422 332279 3478 332288
rect 3436 331375 3464 332279
rect 3422 331366 3478 331375
rect 3422 331301 3478 331310
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324465 580212 325207
rect 580170 324456 580226 324465
rect 580170 324391 580226 324400
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 318321 3464 319223
rect 3422 318312 3478 318321
rect 3422 318247 3478 318256
rect 579618 312080 579674 312089
rect 579618 312015 579674 312024
rect 579526 311128 579582 311137
rect 579632 311114 579660 312015
rect 579582 311086 579660 311114
rect 579526 311063 579582 311072
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 3436 305145 3464 306167
rect 3422 305136 3478 305145
rect 3422 305071 3478 305080
rect 579618 298752 579674 298761
rect 579618 298687 579674 298696
rect 579526 297800 579582 297809
rect 579632 297786 579660 298687
rect 579582 297758 579660 297786
rect 579526 297735 579582 297744
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3436 292091 3464 293111
rect 3422 292082 3478 292091
rect 3422 292017 3478 292026
rect 580170 285424 580226 285433
rect 580170 285359 580226 285368
rect 580184 284481 580212 285359
rect 580170 284472 580226 284481
rect 580170 284407 580226 284416
rect 3422 280120 3478 280129
rect 3422 280055 3478 280064
rect 3436 279037 3464 280055
rect 3422 279028 3478 279037
rect 3422 278963 3478 278972
rect 579618 272232 579674 272241
rect 579618 272167 579674 272176
rect 579526 271144 579582 271153
rect 579632 271130 579660 272167
rect 579582 271102 579660 271130
rect 579526 271079 579582 271088
rect 3422 267200 3478 267209
rect 3422 267135 3478 267144
rect 3436 265983 3464 267135
rect 3422 265974 3478 265983
rect 3422 265909 3478 265918
rect 580906 258904 580962 258913
rect 580906 258839 580962 258848
rect 580920 257854 580948 258839
rect 578884 257848 578936 257854
rect 578884 257790 578936 257796
rect 580908 257848 580960 257854
rect 580908 257790 580960 257796
rect 578896 257689 578924 257790
rect 578882 257680 578938 257689
rect 578882 257615 578938 257624
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3436 252807 3464 254079
rect 3422 252798 3478 252807
rect 3422 252733 3478 252742
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 244497 580212 245511
rect 580170 244488 580226 244497
rect 580170 244423 580226 244432
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3436 239753 3464 241023
rect 3422 239744 3478 239753
rect 3422 239679 3478 239688
rect 579618 232384 579674 232393
rect 579618 232319 579674 232328
rect 579526 231160 579582 231169
rect 579632 231146 579660 232319
rect 579582 231118 579660 231146
rect 579526 231095 579582 231104
rect 3422 228032 3478 228041
rect 3422 227967 3478 227976
rect 3436 226699 3464 227967
rect 3422 226690 3478 226699
rect 3422 226625 3478 226634
rect 579618 219056 579674 219065
rect 579618 218991 579674 219000
rect 579526 217696 579582 217705
rect 579632 217682 579660 218991
rect 579582 217654 579660 217682
rect 579526 217631 579582 217640
rect 3422 214976 3478 214985
rect 3422 214911 3478 214920
rect 3436 213523 3464 214911
rect 3422 213514 3478 213523
rect 3422 213449 3478 213458
rect 579618 205728 579674 205737
rect 579618 205663 579674 205672
rect 579526 204368 579582 204377
rect 579632 204354 579660 205663
rect 579582 204326 579660 204354
rect 579526 204303 579582 204312
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3436 200469 3464 201855
rect 3422 200460 3478 200469
rect 3422 200395 3478 200404
rect 579618 192536 579674 192545
rect 579618 192471 579674 192480
rect 579526 191040 579582 191049
rect 579632 191026 579660 192471
rect 579582 190998 579660 191026
rect 579526 190975 579582 190984
rect 3606 188864 3662 188873
rect 3606 188799 3662 188808
rect 3620 187415 3648 188799
rect 3606 187406 3662 187415
rect 3606 187341 3662 187350
rect 579618 179208 579674 179217
rect 579618 179143 579674 179152
rect 579526 177712 579582 177721
rect 579632 177698 579660 179143
rect 579582 177670 579660 177698
rect 579526 177647 579582 177656
rect 3422 175944 3478 175953
rect 3422 175879 3478 175888
rect 3436 174239 3464 175879
rect 3422 174230 3478 174239
rect 3422 174165 3478 174174
rect 579618 165880 579674 165889
rect 579618 165815 579674 165824
rect 579526 164384 579582 164393
rect 579632 164370 579660 165815
rect 579582 164342 579660 164370
rect 579526 164319 579582 164328
rect 2134 162888 2190 162897
rect 2134 162823 2190 162832
rect 2148 161129 2176 162823
rect 2134 161120 2190 161129
rect 2134 161055 2190 161064
rect 580906 152688 580962 152697
rect 580906 152623 580962 152632
rect 580920 151502 580948 152623
rect 578516 151496 578568 151502
rect 578516 151438 578568 151444
rect 580908 151496 580960 151502
rect 580908 151438 580960 151444
rect 578528 151065 578556 151438
rect 578514 151056 578570 151065
rect 578514 150991 578570 151000
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3436 148131 3464 149767
rect 3422 148122 3478 148131
rect 3422 148057 3478 148066
rect 579618 139360 579674 139369
rect 579618 139295 579674 139304
rect 579526 137592 579582 137601
rect 579632 137578 579660 139295
rect 579582 137550 579660 137578
rect 579526 137527 579582 137536
rect 2134 136776 2190 136785
rect 2134 136711 2190 136720
rect 2148 135017 2176 136711
rect 2134 135008 2190 135017
rect 2134 134943 2190 134952
rect 579618 126032 579674 126041
rect 579618 125967 579674 125976
rect 579526 124400 579582 124409
rect 579632 124386 579660 125967
rect 579582 124358 579660 124386
rect 579526 124335 579582 124344
rect 3422 123720 3478 123729
rect 3422 123655 3478 123664
rect 3436 121901 3464 123655
rect 3422 121892 3478 121901
rect 3422 121827 3478 121836
rect 579618 112840 579674 112849
rect 579618 112775 579674 112784
rect 579526 110936 579582 110945
rect 579632 110922 579660 112775
rect 579582 110894 579660 110922
rect 579526 110871 579582 110880
rect 2134 110664 2190 110673
rect 2134 110599 2190 110608
rect 2148 108905 2176 110599
rect 2134 108896 2190 108905
rect 2134 108831 2190 108840
rect 579618 99512 579674 99521
rect 579618 99447 579674 99456
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 579526 97608 579582 97617
rect 579632 97594 579660 99447
rect 579582 97566 579660 97594
rect 579526 97543 579582 97552
rect 3436 95793 3464 97543
rect 3422 95784 3478 95793
rect 3422 95719 3478 95728
rect 579618 86184 579674 86193
rect 579618 86119 579674 86128
rect 2134 84688 2190 84697
rect 2134 84623 2190 84632
rect 2148 82657 2176 84623
rect 579526 84280 579582 84289
rect 579632 84266 579660 86119
rect 579582 84238 579660 84266
rect 579526 84215 579582 84224
rect 2134 82648 2190 82657
rect 2134 82583 2190 82592
rect 579618 72992 579674 73001
rect 579618 72927 579674 72936
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3436 69563 3464 71567
rect 579526 70952 579582 70961
rect 579632 70938 579660 72927
rect 579582 70910 579660 70938
rect 579526 70887 579582 70896
rect 3422 69554 3478 69563
rect 3422 69489 3478 69498
rect 579618 59664 579674 59673
rect 579618 59599 579674 59608
rect 2134 58576 2190 58585
rect 2134 58511 2190 58520
rect 2148 56545 2176 58511
rect 579526 57624 579582 57633
rect 579632 57610 579660 59599
rect 579582 57582 579660 57610
rect 579526 57559 579582 57568
rect 2134 56536 2190 56545
rect 2134 56471 2190 56480
rect 579986 46336 580042 46345
rect 579986 46271 580042 46280
rect 3422 45520 3478 45529
rect 3422 45455 3478 45464
rect 3436 43333 3464 45455
rect 580000 45014 580028 46271
rect 578332 45008 578384 45014
rect 578332 44950 578384 44956
rect 579988 45008 580040 45014
rect 579988 44950 580040 44956
rect 578344 44305 578372 44950
rect 578330 44296 578386 44305
rect 578330 44231 578386 44240
rect 3422 43324 3478 43333
rect 3422 43259 3478 43268
rect 579618 33144 579674 33153
rect 579618 33079 579674 33088
rect 2134 32464 2190 32473
rect 2134 32399 2190 32408
rect 2148 30297 2176 32399
rect 579526 30968 579582 30977
rect 579632 30954 579660 33079
rect 579582 30926 579660 30954
rect 579526 30903 579582 30912
rect 2134 30288 2190 30297
rect 2134 30223 2190 30232
rect 579618 19816 579674 19825
rect 579618 19751 579674 19760
rect 2042 19408 2098 19417
rect 2042 19343 2098 19352
rect 2056 17241 2084 19343
rect 579526 17640 579582 17649
rect 579632 17626 579660 19751
rect 579582 17598 579660 17626
rect 579526 17575 579582 17584
rect 2042 17232 2098 17241
rect 2042 17167 2098 17176
rect 579618 6624 579674 6633
rect 579618 6559 579674 6568
rect 2778 6488 2834 6497
rect 2778 6423 2834 6432
rect 2792 4185 2820 6423
rect 579632 5574 579660 6559
rect 576860 5568 576912 5574
rect 576860 5510 576912 5516
rect 579620 5568 579672 5574
rect 579620 5510 579672 5516
rect 2778 4176 2834 4185
rect 2778 4111 2834 4120
rect 576766 4176 576822 4185
rect 576872 4162 576900 5510
rect 576822 4134 576900 4162
rect 576766 4111 576822 4120
rect 1676 3868 1728 3874
rect 1676 3810 1728 3816
rect 572 3800 624 3806
rect 572 3742 624 3748
rect 584 480 612 3742
rect 1688 480 1716 3810
rect 4124 3806 4152 4012
rect 5228 3874 5256 4012
rect 5216 3868 5268 3874
rect 5216 3810 5268 3816
rect 4112 3800 4164 3806
rect 6424 3754 6452 4012
rect 7528 3754 7556 4012
rect 4112 3742 4164 3748
rect 6380 3726 6452 3754
rect 7484 3726 7556 3754
rect 7656 3800 7708 3806
rect 8724 3754 8752 4012
rect 9920 3754 9948 4012
rect 11024 3806 11052 4012
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 7656 3742 7708 3748
rect 4068 2848 4120 2854
rect 4068 2790 4120 2796
rect 3240 1352 3292 1358
rect 3240 1294 3292 1300
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 354 2954 480
rect 3252 354 3280 1294
rect 4080 480 4108 2790
rect 6380 1358 6408 3726
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6368 1352 6420 1358
rect 6368 1294 6420 1300
rect 5632 1148 5684 1154
rect 5632 1090 5684 1096
rect 2842 326 3280 354
rect 2842 -960 2954 326
rect 4038 -960 4150 480
rect 5234 354 5346 480
rect 5644 354 5672 1090
rect 6472 480 6500 2994
rect 7484 2854 7512 3726
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7668 480 7696 3742
rect 8680 3726 8752 3754
rect 9876 3726 9948 3754
rect 11012 3800 11064 3806
rect 11012 3742 11064 3748
rect 8680 1154 8708 3726
rect 9876 3058 9904 3726
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 8668 1148 8720 1154
rect 8668 1090 8720 1096
rect 8760 944 8812 950
rect 8760 886 8812 892
rect 8772 480 8800 886
rect 9968 480 9996 2790
rect 11164 480 11192 3878
rect 12220 3754 12248 4012
rect 12176 3726 12248 3754
rect 12348 3800 12400 3806
rect 13324 3754 13352 4012
rect 14520 3942 14548 4012
rect 14508 3936 14560 3942
rect 14508 3878 14560 3884
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 13544 3868 13596 3874
rect 13544 3810 13596 3816
rect 12348 3742 12400 3748
rect 12176 950 12204 3726
rect 12164 944 12216 950
rect 12164 886 12216 892
rect 12360 480 12388 3742
rect 13280 3726 13352 3754
rect 13280 2854 13308 3726
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 13556 480 13584 3810
rect 14752 480 14780 3878
rect 15716 3806 15744 4012
rect 16820 3874 16848 4012
rect 18016 3942 18044 4012
rect 18004 3936 18056 3942
rect 18004 3878 18056 3884
rect 16808 3868 16860 3874
rect 16808 3810 16860 3816
rect 19120 3806 19148 4012
rect 19432 3868 19484 3874
rect 19432 3810 19484 3816
rect 15704 3800 15756 3806
rect 15704 3742 15756 3748
rect 15936 3800 15988 3806
rect 15936 3742 15988 3748
rect 19108 3800 19160 3806
rect 19108 3742 19160 3748
rect 15948 480 15976 3742
rect 18236 2916 18288 2922
rect 18236 2858 18288 2864
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 17052 480 17080 2790
rect 18248 480 18276 2858
rect 19444 480 19472 3810
rect 20316 3754 20344 4012
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20272 3726 20344 3754
rect 20272 2854 20300 3726
rect 20260 2848 20312 2854
rect 20260 2790 20312 2796
rect 20640 480 20668 3878
rect 21512 3754 21540 4012
rect 22616 3874 22644 4012
rect 23812 3942 23840 4012
rect 23800 3936 23852 3942
rect 23800 3878 23852 3884
rect 24216 3936 24268 3942
rect 24216 3878 24268 3884
rect 22604 3868 22656 3874
rect 22604 3810 22656 3816
rect 23020 3868 23072 3874
rect 23020 3810 23072 3816
rect 21468 3726 21540 3754
rect 21824 3800 21876 3806
rect 21824 3742 21876 3748
rect 21468 2922 21496 3726
rect 21456 2916 21508 2922
rect 21456 2858 21508 2864
rect 21836 480 21864 3742
rect 23032 480 23060 3810
rect 24228 480 24256 3878
rect 24916 3806 24944 4012
rect 26112 3874 26140 4012
rect 27308 3942 27336 4012
rect 27296 3936 27348 3942
rect 27296 3878 27348 3884
rect 27712 3936 27764 3942
rect 27712 3878 27764 3884
rect 26100 3868 26152 3874
rect 26100 3810 26152 3816
rect 26516 3868 26568 3874
rect 26516 3810 26568 3816
rect 24904 3800 24956 3806
rect 24904 3742 24956 3748
rect 25320 3800 25372 3806
rect 25320 3742 25372 3748
rect 25332 480 25360 3742
rect 26528 480 26556 3810
rect 27724 480 27752 3878
rect 28412 3806 28440 4012
rect 29608 3874 29636 4012
rect 30712 3942 30740 4012
rect 30700 3936 30752 3942
rect 30700 3878 30752 3884
rect 29596 3868 29648 3874
rect 29596 3810 29648 3816
rect 30104 3868 30156 3874
rect 30104 3810 30156 3816
rect 28400 3800 28452 3806
rect 28400 3742 28452 3748
rect 28908 2848 28960 2854
rect 28908 2790 28960 2796
rect 28920 480 28948 2790
rect 30116 480 30144 3810
rect 31300 3800 31352 3806
rect 31908 3754 31936 4012
rect 32404 3936 32456 3942
rect 32404 3878 32456 3884
rect 31300 3742 31352 3748
rect 31312 480 31340 3742
rect 31864 3726 31936 3754
rect 31864 2854 31892 3726
rect 31852 2848 31904 2854
rect 31852 2790 31904 2796
rect 32416 480 32444 3878
rect 33104 3874 33132 4012
rect 33092 3868 33144 3874
rect 33092 3810 33144 3816
rect 33600 3868 33652 3874
rect 33600 3810 33652 3816
rect 33612 480 33640 3810
rect 34208 3806 34236 4012
rect 35404 3942 35432 4012
rect 35392 3936 35444 3942
rect 35392 3878 35444 3884
rect 36600 3874 36628 4012
rect 36588 3868 36640 3874
rect 36588 3810 36640 3816
rect 37188 3868 37240 3874
rect 37188 3810 37240 3816
rect 34196 3800 34248 3806
rect 34196 3742 34248 3748
rect 34796 3800 34848 3806
rect 34796 3742 34848 3748
rect 34808 480 34836 3742
rect 35992 2848 36044 2854
rect 35992 2790 36044 2796
rect 36004 480 36032 2790
rect 37200 480 37228 3810
rect 37704 3806 37732 4012
rect 38384 3936 38436 3942
rect 38384 3878 38436 3884
rect 37692 3800 37744 3806
rect 37692 3742 37744 3748
rect 38396 480 38424 3878
rect 38900 3754 38928 4012
rect 40004 3874 40032 4012
rect 41200 3942 41228 4012
rect 41188 3936 41240 3942
rect 41188 3878 41240 3884
rect 39992 3868 40044 3874
rect 39992 3810 40044 3816
rect 41880 3868 41932 3874
rect 41880 3810 41932 3816
rect 38856 3726 38928 3754
rect 40684 3800 40736 3806
rect 40684 3742 40736 3748
rect 38856 2854 38884 3726
rect 38844 2848 38896 2854
rect 38844 2790 38896 2796
rect 39580 2848 39632 2854
rect 39580 2790 39632 2796
rect 39592 480 39620 2790
rect 40696 480 40724 3742
rect 41892 480 41920 3810
rect 42396 3754 42424 4012
rect 43076 3936 43128 3942
rect 43076 3878 43128 3884
rect 42352 3726 42424 3754
rect 42352 2854 42380 3726
rect 42340 2848 42392 2854
rect 42340 2790 42392 2796
rect 43088 480 43116 3878
rect 43500 3806 43528 4012
rect 44696 3874 44724 4012
rect 45800 3942 45828 4012
rect 45788 3936 45840 3942
rect 45788 3878 45840 3884
rect 46664 3936 46716 3942
rect 46664 3878 46716 3884
rect 44684 3868 44736 3874
rect 44684 3810 44736 3816
rect 45468 3868 45520 3874
rect 45468 3810 45520 3816
rect 43488 3800 43540 3806
rect 43488 3742 43540 3748
rect 44272 3800 44324 3806
rect 44272 3742 44324 3748
rect 44284 480 44312 3742
rect 45480 480 45508 3810
rect 46676 480 46704 3878
rect 46996 3806 47024 4012
rect 48192 3874 48220 4012
rect 49296 3942 49324 4012
rect 49284 3936 49336 3942
rect 49284 3878 49336 3884
rect 50160 3936 50212 3942
rect 50160 3878 50212 3884
rect 48180 3868 48232 3874
rect 48180 3810 48232 3816
rect 48964 3868 49016 3874
rect 48964 3810 49016 3816
rect 46984 3800 47036 3806
rect 46984 3742 47036 3748
rect 47860 3800 47912 3806
rect 47860 3742 47912 3748
rect 47872 480 47900 3742
rect 48976 480 49004 3810
rect 50172 480 50200 3878
rect 50492 3806 50520 4012
rect 51596 3874 51624 4012
rect 52792 3942 52820 4012
rect 52780 3936 52832 3942
rect 52780 3878 52832 3884
rect 51584 3868 51636 3874
rect 51584 3810 51636 3816
rect 53748 3868 53800 3874
rect 53748 3810 53800 3816
rect 50480 3800 50532 3806
rect 50480 3742 50532 3748
rect 51356 3800 51408 3806
rect 51356 3742 51408 3748
rect 51368 480 51396 3742
rect 52552 740 52604 746
rect 52552 682 52604 688
rect 52564 480 52592 682
rect 53760 480 53788 3810
rect 53988 3806 54016 4012
rect 53976 3800 54028 3806
rect 53976 3742 54028 3748
rect 54944 3800 54996 3806
rect 55092 3754 55120 4012
rect 56048 3936 56100 3942
rect 56048 3878 56100 3884
rect 54944 3742 54996 3748
rect 54956 480 54984 3742
rect 55048 3726 55120 3754
rect 55048 746 55076 3726
rect 55036 740 55088 746
rect 55036 682 55088 688
rect 56060 480 56088 3878
rect 56288 3874 56316 4012
rect 56276 3868 56328 3874
rect 56276 3810 56328 3816
rect 57244 3868 57296 3874
rect 57244 3810 57296 3816
rect 57256 480 57284 3810
rect 57392 3806 57420 4012
rect 58588 3942 58616 4012
rect 58576 3936 58628 3942
rect 58576 3878 58628 3884
rect 59784 3874 59812 4012
rect 59772 3868 59824 3874
rect 59772 3810 59824 3816
rect 60888 3806 60916 4012
rect 62084 3890 62112 4012
rect 61948 3862 62112 3890
rect 57380 3800 57432 3806
rect 57380 3742 57432 3748
rect 58440 3800 58492 3806
rect 58440 3742 58492 3748
rect 60876 3800 60928 3806
rect 60876 3742 60928 3748
rect 58452 480 58480 3742
rect 60832 1352 60884 1358
rect 60832 1294 60884 1300
rect 59636 740 59688 746
rect 59636 682 59688 688
rect 59648 480 59676 682
rect 60844 480 60872 1294
rect 61948 746 61976 3862
rect 63280 3754 63308 4012
rect 64384 3890 64412 4012
rect 64384 3862 64460 3890
rect 64328 3800 64380 3806
rect 63280 3726 63356 3754
rect 64328 3742 64380 3748
rect 63224 3052 63276 3058
rect 63224 2994 63276 3000
rect 62028 2848 62080 2854
rect 62028 2790 62080 2796
rect 61936 740 61988 746
rect 61936 682 61988 688
rect 62040 480 62068 2790
rect 63236 480 63264 2994
rect 63328 1358 63356 3726
rect 63316 1352 63368 1358
rect 63316 1294 63368 1300
rect 64340 480 64368 3742
rect 64432 2854 64460 3862
rect 65580 3754 65608 4012
rect 66684 3806 66712 4012
rect 65536 3726 65608 3754
rect 66672 3800 66724 3806
rect 66672 3742 66724 3748
rect 67088 3800 67140 3806
rect 67880 3754 67908 4012
rect 69076 3806 69104 4012
rect 67088 3742 67140 3748
rect 65536 3058 65564 3726
rect 65524 3052 65576 3058
rect 65524 2994 65576 3000
rect 64420 2848 64472 2854
rect 64420 2790 64472 2796
rect 65524 2848 65576 2854
rect 65524 2790 65576 2796
rect 65536 480 65564 2790
rect 5234 326 5672 354
rect 5234 -960 5346 326
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 354 66802 480
rect 67100 354 67128 3742
rect 67836 3726 67908 3754
rect 69064 3800 69116 3806
rect 70180 3754 70208 4012
rect 69064 3742 69116 3748
rect 70136 3726 70208 3754
rect 70308 3800 70360 3806
rect 71376 3754 71404 4012
rect 71504 3868 71556 3874
rect 71504 3810 71556 3816
rect 70308 3742 70360 3748
rect 67836 2854 67864 3726
rect 67824 2848 67876 2854
rect 67824 2790 67876 2796
rect 70136 1358 70164 3726
rect 67916 1352 67968 1358
rect 67916 1294 67968 1300
rect 70124 1352 70176 1358
rect 70124 1294 70176 1300
rect 67928 480 67956 1294
rect 69112 604 69164 610
rect 69112 546 69164 552
rect 69124 480 69152 546
rect 70320 480 70348 3742
rect 71332 3726 71404 3754
rect 71332 610 71360 3726
rect 71320 604 71372 610
rect 71320 546 71372 552
rect 71516 480 71544 3810
rect 72480 3806 72508 4012
rect 72608 3936 72660 3942
rect 72608 3878 72660 3884
rect 72468 3800 72520 3806
rect 72468 3742 72520 3748
rect 72620 480 72648 3878
rect 73676 3874 73704 4012
rect 74872 3942 74900 4012
rect 74860 3936 74912 3942
rect 74860 3878 74912 3884
rect 73664 3868 73716 3874
rect 73664 3810 73716 3816
rect 75976 3806 76004 4012
rect 73804 3800 73856 3806
rect 73804 3742 73856 3748
rect 75964 3800 76016 3806
rect 77172 3754 77200 4012
rect 78276 3754 78304 4012
rect 78588 3868 78640 3874
rect 78588 3810 78640 3816
rect 75964 3742 76016 3748
rect 73816 480 73844 3742
rect 77128 3726 77200 3754
rect 78232 3726 78304 3754
rect 76196 1352 76248 1358
rect 76196 1294 76248 1300
rect 75000 1284 75052 1290
rect 75000 1226 75052 1232
rect 75012 480 75040 1226
rect 76208 480 76236 1294
rect 77128 1290 77156 3726
rect 78232 1358 78260 3726
rect 78220 1352 78272 1358
rect 78220 1294 78272 1300
rect 77116 1284 77168 1290
rect 77116 1226 77168 1232
rect 77392 1284 77444 1290
rect 77392 1226 77444 1232
rect 77404 480 77432 1226
rect 78600 480 78628 3810
rect 79472 3754 79500 4012
rect 80668 3874 80696 4012
rect 80656 3868 80708 3874
rect 80656 3810 80708 3816
rect 80888 3868 80940 3874
rect 80888 3810 80940 3816
rect 79428 3726 79500 3754
rect 79692 3800 79744 3806
rect 79692 3742 79744 3748
rect 79428 1290 79456 3726
rect 79416 1284 79468 1290
rect 79416 1226 79468 1232
rect 79704 480 79732 3742
rect 80900 480 80928 3810
rect 81772 3806 81800 4012
rect 82968 3874 82996 4012
rect 82956 3868 83008 3874
rect 82956 3810 83008 3816
rect 81760 3800 81812 3806
rect 84072 3754 84100 4012
rect 85268 3754 85296 4012
rect 86464 3754 86492 4012
rect 81760 3742 81812 3748
rect 84028 3726 84100 3754
rect 85224 3726 85296 3754
rect 86420 3726 86492 3754
rect 86868 3800 86920 3806
rect 87568 3754 87596 4012
rect 87972 3868 88024 3874
rect 87972 3810 88024 3816
rect 86868 3742 86920 3748
rect 83280 1352 83332 1358
rect 83280 1294 83332 1300
rect 82084 1284 82136 1290
rect 82084 1226 82136 1232
rect 82096 480 82124 1226
rect 83292 480 83320 1294
rect 84028 1290 84056 3726
rect 85224 1358 85252 3726
rect 85212 1352 85264 1358
rect 85212 1294 85264 1300
rect 85672 1352 85724 1358
rect 85672 1294 85724 1300
rect 84016 1284 84068 1290
rect 84016 1226 84068 1232
rect 84476 1284 84528 1290
rect 84476 1226 84528 1232
rect 84488 480 84516 1226
rect 85684 480 85712 1294
rect 86420 1290 86448 3726
rect 86408 1284 86460 1290
rect 86408 1226 86460 1232
rect 86880 480 86908 3742
rect 87524 3726 87596 3754
rect 87524 1358 87552 3726
rect 87512 1352 87564 1358
rect 87512 1294 87564 1300
rect 87984 480 88012 3810
rect 88764 3806 88792 4012
rect 89960 3874 89988 4012
rect 89948 3868 90000 3874
rect 89948 3810 90000 3816
rect 88752 3800 88804 3806
rect 91064 3754 91092 4012
rect 92260 3754 92288 4012
rect 93364 3754 93392 4012
rect 94560 3754 94588 4012
rect 88752 3742 88804 3748
rect 91020 3726 91092 3754
rect 92216 3726 92288 3754
rect 93320 3726 93392 3754
rect 94516 3726 94588 3754
rect 95148 3800 95200 3806
rect 95756 3754 95784 4012
rect 96252 3868 96304 3874
rect 96252 3810 96304 3816
rect 95148 3742 95200 3748
rect 91020 1358 91048 3726
rect 89168 1352 89220 1358
rect 89168 1294 89220 1300
rect 91008 1352 91060 1358
rect 91008 1294 91060 1300
rect 91560 1352 91612 1358
rect 91560 1294 91612 1300
rect 89180 480 89208 1294
rect 90364 1284 90416 1290
rect 90364 1226 90416 1232
rect 90376 480 90404 1226
rect 91572 480 91600 1294
rect 92216 1290 92244 3726
rect 93320 1358 93348 3726
rect 93308 1352 93360 1358
rect 93308 1294 93360 1300
rect 93952 1352 94004 1358
rect 93952 1294 94004 1300
rect 92204 1284 92256 1290
rect 92204 1226 92256 1232
rect 92756 1284 92808 1290
rect 92756 1226 92808 1232
rect 92768 480 92796 1226
rect 93964 480 93992 1294
rect 94516 1290 94544 3726
rect 94504 1284 94556 1290
rect 94504 1226 94556 1232
rect 95160 480 95188 3742
rect 95712 3726 95784 3754
rect 95712 1358 95740 3726
rect 95700 1352 95752 1358
rect 95700 1294 95752 1300
rect 96264 480 96292 3810
rect 96860 3806 96888 4012
rect 98056 3874 98084 4012
rect 98044 3868 98096 3874
rect 98044 3810 98096 3816
rect 96848 3800 96900 3806
rect 99160 3754 99188 4012
rect 100356 3754 100384 4012
rect 101552 3754 101580 4012
rect 102656 3754 102684 4012
rect 96848 3742 96900 3748
rect 99116 3726 99188 3754
rect 100312 3726 100384 3754
rect 101508 3726 101580 3754
rect 102612 3726 102684 3754
rect 103336 3800 103388 3806
rect 103852 3754 103880 4012
rect 104956 3806 104984 4012
rect 103336 3742 103388 3748
rect 99116 1358 99144 3726
rect 97448 1352 97500 1358
rect 97448 1294 97500 1300
rect 99104 1352 99156 1358
rect 99104 1294 99156 1300
rect 97460 480 97488 1294
rect 100312 1290 100340 3726
rect 101036 1352 101088 1358
rect 101036 1294 101088 1300
rect 98644 1284 98696 1290
rect 98644 1226 98696 1232
rect 100300 1284 100352 1290
rect 100300 1226 100352 1232
rect 98656 480 98684 1226
rect 99840 1216 99892 1222
rect 99840 1158 99892 1164
rect 99852 480 99880 1158
rect 101048 480 101076 1294
rect 101508 1222 101536 3726
rect 102612 1358 102640 3726
rect 102600 1352 102652 1358
rect 102600 1294 102652 1300
rect 102232 1284 102284 1290
rect 102232 1226 102284 1232
rect 101496 1216 101548 1222
rect 101496 1158 101548 1164
rect 102244 480 102272 1226
rect 103348 480 103376 3742
rect 103808 3726 103880 3754
rect 104944 3800 104996 3806
rect 106152 3754 106180 4012
rect 107348 3754 107376 4012
rect 108452 3754 108480 4012
rect 109648 3754 109676 4012
rect 110752 3754 110780 4012
rect 111948 3754 111976 4012
rect 113144 3754 113172 4012
rect 114248 3754 114276 4012
rect 115444 3754 115472 4012
rect 116640 3754 116668 4012
rect 117744 3754 117772 4012
rect 118940 3754 118968 4012
rect 120044 3754 120072 4012
rect 121240 3754 121268 4012
rect 122436 3754 122464 4012
rect 123540 3754 123568 4012
rect 104944 3742 104996 3748
rect 106108 3726 106180 3754
rect 107304 3726 107376 3754
rect 108408 3726 108480 3754
rect 109604 3726 109676 3754
rect 110708 3726 110780 3754
rect 111904 3726 111976 3754
rect 113100 3726 113172 3754
rect 114204 3726 114276 3754
rect 115400 3726 115472 3754
rect 116596 3726 116668 3754
rect 117700 3726 117772 3754
rect 118896 3726 118968 3754
rect 119264 3726 120072 3754
rect 121196 3726 121268 3754
rect 122392 3726 122464 3754
rect 123496 3726 123568 3754
rect 124736 3754 124764 4012
rect 125840 3754 125868 4012
rect 127036 3754 127064 4012
rect 128232 3754 128260 4012
rect 129336 3754 129364 4012
rect 130532 3754 130560 4012
rect 131636 3754 131664 4012
rect 132832 3754 132860 4012
rect 134028 3754 134056 4012
rect 135132 3754 135160 4012
rect 136328 3754 136356 4012
rect 137432 3754 137460 4012
rect 138628 3754 138656 4012
rect 139824 3754 139852 4012
rect 140928 3754 140956 4012
rect 142124 3754 142152 4012
rect 143320 3754 143348 4012
rect 144424 3754 144452 4012
rect 145620 3754 145648 4012
rect 146724 3754 146752 4012
rect 147920 3754 147948 4012
rect 149116 3754 149144 4012
rect 150220 3754 150248 4012
rect 151416 3754 151444 4012
rect 152520 3754 152548 4012
rect 153716 3754 153744 4012
rect 154912 3754 154940 4012
rect 156016 3754 156044 4012
rect 157212 3754 157240 4012
rect 158316 3754 158344 4012
rect 159512 3754 159540 4012
rect 160708 3754 160736 4012
rect 161812 3754 161840 4012
rect 163008 3754 163036 4012
rect 164112 3754 164140 4012
rect 165308 3754 165336 4012
rect 166504 3754 166532 4012
rect 167608 3754 167636 4012
rect 168804 3754 168832 4012
rect 170000 3754 170028 4012
rect 171104 3754 171132 4012
rect 172300 3754 172328 4012
rect 173404 3754 173432 4012
rect 174600 3754 174628 4012
rect 175796 3754 175824 4012
rect 176900 3754 176928 4012
rect 178096 3754 178124 4012
rect 179200 3754 179228 4012
rect 124736 3726 124812 3754
rect 103808 1290 103836 3726
rect 106108 1358 106136 3726
rect 104532 1352 104584 1358
rect 104532 1294 104584 1300
rect 106096 1352 106148 1358
rect 106096 1294 106148 1300
rect 106924 1352 106976 1358
rect 106924 1294 106976 1300
rect 103796 1284 103848 1290
rect 103796 1226 103848 1232
rect 104544 480 104572 1294
rect 105728 740 105780 746
rect 105728 682 105780 688
rect 105740 480 105768 682
rect 106936 480 106964 1294
rect 107304 746 107332 3726
rect 108408 1358 108436 3726
rect 108396 1352 108448 1358
rect 108396 1294 108448 1300
rect 109316 1352 109368 1358
rect 109316 1294 109368 1300
rect 108120 1284 108172 1290
rect 108120 1226 108172 1232
rect 107292 740 107344 746
rect 107292 682 107344 688
rect 108132 480 108160 1226
rect 109328 480 109356 1294
rect 109604 1290 109632 3726
rect 110708 1358 110736 3726
rect 110696 1352 110748 1358
rect 110696 1294 110748 1300
rect 111904 1290 111932 3726
rect 112812 1352 112864 1358
rect 112812 1294 112864 1300
rect 109592 1284 109644 1290
rect 109592 1226 109644 1232
rect 110512 1284 110564 1290
rect 110512 1226 110564 1232
rect 111892 1284 111944 1290
rect 111892 1226 111944 1232
rect 110524 480 110552 1226
rect 111616 1148 111668 1154
rect 111616 1090 111668 1096
rect 111628 480 111656 1090
rect 112824 480 112852 1294
rect 113100 1154 113128 3726
rect 114204 1358 114232 3726
rect 114192 1352 114244 1358
rect 114192 1294 114244 1300
rect 115204 1284 115256 1290
rect 115204 1226 115256 1232
rect 114008 1216 114060 1222
rect 114008 1158 114060 1164
rect 113088 1148 113140 1154
rect 113088 1090 113140 1096
rect 114020 480 114048 1158
rect 115216 480 115244 1226
rect 115400 1222 115428 3726
rect 116400 1352 116452 1358
rect 116400 1294 116452 1300
rect 115388 1216 115440 1222
rect 115388 1158 115440 1164
rect 116412 480 116440 1294
rect 116596 1290 116624 3726
rect 117700 1358 117728 3726
rect 117688 1352 117740 1358
rect 117688 1294 117740 1300
rect 118896 1290 118924 3726
rect 116584 1284 116636 1290
rect 116584 1226 116636 1232
rect 117596 1284 117648 1290
rect 117596 1226 117648 1232
rect 118884 1284 118936 1290
rect 118884 1226 118936 1232
rect 117608 480 117636 1226
rect 66690 326 67128 354
rect 66690 -960 66802 326
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 354 118874 480
rect 119264 354 119292 3726
rect 121196 1358 121224 3726
rect 119896 1352 119948 1358
rect 119896 1294 119948 1300
rect 121184 1352 121236 1358
rect 121184 1294 121236 1300
rect 119908 480 119936 1294
rect 122288 1284 122340 1290
rect 122288 1226 122340 1232
rect 121092 944 121144 950
rect 121092 886 121144 892
rect 121104 480 121132 886
rect 122300 480 122328 1226
rect 122392 950 122420 3726
rect 123496 1290 123524 3726
rect 123484 1284 123536 1290
rect 123484 1226 123536 1232
rect 124680 1284 124732 1290
rect 124680 1226 124732 1232
rect 123484 1148 123536 1154
rect 123484 1090 123536 1096
rect 122380 944 122432 950
rect 122380 886 122432 892
rect 123496 480 123524 1090
rect 124692 480 124720 1226
rect 124784 1154 124812 3726
rect 125796 3726 125868 3754
rect 126992 3726 127064 3754
rect 127176 3726 128260 3754
rect 129292 3726 129364 3754
rect 130488 3726 130560 3754
rect 131592 3726 131664 3754
rect 132788 3726 132860 3754
rect 133984 3726 134056 3754
rect 134168 3726 135160 3754
rect 135272 3726 136356 3754
rect 137388 3726 137460 3754
rect 138584 3726 138656 3754
rect 139780 3726 139852 3754
rect 140884 3726 140956 3754
rect 141712 3726 142152 3754
rect 142448 3726 143348 3754
rect 143552 3726 144452 3754
rect 145576 3726 145648 3754
rect 146680 3726 146752 3754
rect 147600 3726 147948 3754
rect 149072 3726 149144 3754
rect 149992 3726 150248 3754
rect 151096 3726 151444 3754
rect 151832 3726 152548 3754
rect 153488 3726 153744 3754
rect 154868 3726 154940 3754
rect 155880 3726 156044 3754
rect 156616 3726 157240 3754
rect 158272 3726 158344 3754
rect 159376 3726 159540 3754
rect 160112 3726 160736 3754
rect 161584 3726 161840 3754
rect 162964 3726 163036 3754
rect 164068 3726 164140 3754
rect 164896 3726 165336 3754
rect 166460 3726 166532 3754
rect 167564 3726 167636 3754
rect 168392 3726 168832 3754
rect 169956 3726 170028 3754
rect 170784 3726 171132 3754
rect 172256 3726 172328 3754
rect 173176 3726 173432 3754
rect 174280 3726 174628 3754
rect 175752 3726 175824 3754
rect 176672 3726 176928 3754
rect 178052 3726 178124 3754
rect 179064 3726 179228 3754
rect 180396 3754 180424 4012
rect 181592 3754 181620 4012
rect 182696 3754 182724 4012
rect 180396 3726 180472 3754
rect 125796 1290 125824 3726
rect 126992 1358 127020 3726
rect 125876 1352 125928 1358
rect 125876 1294 125928 1300
rect 126980 1352 127032 1358
rect 126980 1294 127032 1300
rect 125784 1284 125836 1290
rect 125784 1226 125836 1232
rect 124772 1148 124824 1154
rect 124772 1090 124824 1096
rect 125888 480 125916 1294
rect 127176 1170 127204 3726
rect 129292 1290 129320 3726
rect 130488 1358 130516 3726
rect 131592 1358 131620 3726
rect 132788 1358 132816 3726
rect 133984 1358 134012 3726
rect 129372 1352 129424 1358
rect 129372 1294 129424 1300
rect 130476 1352 130528 1358
rect 130476 1294 130528 1300
rect 130568 1352 130620 1358
rect 130568 1294 130620 1300
rect 131580 1352 131632 1358
rect 131580 1294 131632 1300
rect 131764 1352 131816 1358
rect 131764 1294 131816 1300
rect 132776 1352 132828 1358
rect 132776 1294 132828 1300
rect 132960 1352 133012 1358
rect 132960 1294 133012 1300
rect 133972 1352 134024 1358
rect 133972 1294 134024 1300
rect 128176 1284 128228 1290
rect 128176 1226 128228 1232
rect 129280 1284 129332 1290
rect 129280 1226 129332 1232
rect 126992 1142 127204 1170
rect 126992 480 127020 1142
rect 128188 480 128216 1226
rect 129384 480 129412 1294
rect 130580 480 130608 1294
rect 131776 480 131804 1294
rect 132972 480 133000 1294
rect 134168 480 134196 3726
rect 135272 480 135300 3726
rect 137388 1290 137416 3726
rect 138584 1358 138612 3726
rect 137652 1352 137704 1358
rect 137652 1294 137704 1300
rect 138572 1352 138624 1358
rect 138572 1294 138624 1300
rect 136456 1284 136508 1290
rect 136456 1226 136508 1232
rect 137376 1284 137428 1290
rect 137376 1226 137428 1232
rect 136468 480 136496 1226
rect 137664 480 137692 1294
rect 139780 1290 139808 3726
rect 140884 1290 140912 3726
rect 138848 1284 138900 1290
rect 138848 1226 138900 1232
rect 139768 1284 139820 1290
rect 139768 1226 139820 1232
rect 140044 1284 140096 1290
rect 140044 1226 140096 1232
rect 140872 1284 140924 1290
rect 140872 1226 140924 1232
rect 138860 480 138888 1226
rect 140056 480 140084 1226
rect 118762 326 119292 354
rect 118762 -960 118874 326
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 354 141322 480
rect 141712 354 141740 3726
rect 142448 480 142476 3726
rect 143552 480 143580 3726
rect 145576 1358 145604 3726
rect 146680 1358 146708 3726
rect 144736 1352 144788 1358
rect 144736 1294 144788 1300
rect 145564 1352 145616 1358
rect 145564 1294 145616 1300
rect 145932 1352 145984 1358
rect 145932 1294 145984 1300
rect 146668 1352 146720 1358
rect 146668 1294 146720 1300
rect 144748 480 144776 1294
rect 145944 480 145972 1294
rect 141210 326 141740 354
rect 141210 -960 141322 326
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 354 147210 480
rect 147600 354 147628 3726
rect 149072 1358 149100 3726
rect 148324 1352 148376 1358
rect 148324 1294 148376 1300
rect 149060 1352 149112 1358
rect 149060 1294 149112 1300
rect 148336 480 148364 1294
rect 147098 326 147628 354
rect 147098 -960 147210 326
rect 148294 -960 148406 480
rect 149490 354 149602 480
rect 149992 354 150020 3726
rect 149490 326 150020 354
rect 150594 354 150706 480
rect 151096 354 151124 3726
rect 151832 480 151860 3726
rect 150594 326 151124 354
rect 149490 -960 149602 326
rect 150594 -960 150706 326
rect 151790 -960 151902 480
rect 152986 354 153098 480
rect 153488 354 153516 3726
rect 154868 1358 154896 3726
rect 154212 1352 154264 1358
rect 154212 1294 154264 1300
rect 154856 1352 154908 1358
rect 154856 1294 154908 1300
rect 154224 480 154252 1294
rect 152986 326 153516 354
rect 152986 -960 153098 326
rect 154182 -960 154294 480
rect 155378 354 155490 480
rect 155880 354 155908 3726
rect 156616 480 156644 3726
rect 155378 326 155908 354
rect 155378 -960 155490 326
rect 156574 -960 156686 480
rect 157770 354 157882 480
rect 158272 354 158300 3726
rect 157770 326 158300 354
rect 158874 354 158986 480
rect 159376 354 159404 3726
rect 160112 480 160140 3726
rect 158874 326 159404 354
rect 157770 -960 157882 326
rect 158874 -960 158986 326
rect 160070 -960 160182 480
rect 161266 354 161378 480
rect 161584 354 161612 3726
rect 162964 1358 162992 3726
rect 162492 1352 162544 1358
rect 162492 1294 162544 1300
rect 162952 1352 163004 1358
rect 162952 1294 163004 1300
rect 162504 480 162532 1294
rect 161266 326 161612 354
rect 161266 -960 161378 326
rect 162462 -960 162574 480
rect 163658 354 163770 480
rect 164068 354 164096 3726
rect 164896 480 164924 3726
rect 163658 326 164096 354
rect 163658 -960 163770 326
rect 164854 -960 164966 480
rect 166050 354 166162 480
rect 166460 354 166488 3726
rect 166050 326 166488 354
rect 167154 354 167266 480
rect 167564 354 167592 3726
rect 168392 480 168420 3726
rect 167154 326 167592 354
rect 166050 -960 166162 326
rect 167154 -960 167266 326
rect 168350 -960 168462 480
rect 169546 354 169658 480
rect 169956 354 169984 3726
rect 170784 480 170812 3726
rect 169546 326 169984 354
rect 169546 -960 169658 326
rect 170742 -960 170854 480
rect 171938 354 172050 480
rect 172256 354 172284 3726
rect 173176 480 173204 3726
rect 174280 480 174308 3726
rect 171938 326 172284 354
rect 171938 -960 172050 326
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 354 175546 480
rect 175752 354 175780 3726
rect 176672 480 176700 3726
rect 175434 326 175780 354
rect 175434 -960 175546 326
rect 176630 -960 176742 480
rect 177826 354 177938 480
rect 178052 354 178080 3726
rect 179064 480 179092 3726
rect 177826 326 178080 354
rect 177826 -960 177938 326
rect 179022 -960 179134 480
rect 180218 218 180330 480
rect 180444 218 180472 3726
rect 181456 3726 181620 3754
rect 182560 3726 182724 3754
rect 183892 3754 183920 4012
rect 184996 3754 185024 4012
rect 186192 3754 186220 4012
rect 187388 3754 187416 4012
rect 183892 3726 183968 3754
rect 181456 480 181484 3726
rect 182560 480 182588 3726
rect 180218 190 180472 218
rect 180218 -960 180330 190
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 218 183826 480
rect 183940 218 183968 3726
rect 184952 3726 185024 3754
rect 186148 3726 186220 3754
rect 187344 3726 187416 3754
rect 188492 3754 188520 4012
rect 189688 3754 189716 4012
rect 190792 3754 190820 4012
rect 191988 3754 192016 4012
rect 193184 3754 193212 4012
rect 194288 3754 194316 4012
rect 195484 3754 195512 4012
rect 188492 3726 188568 3754
rect 189688 3726 189764 3754
rect 190792 3726 190868 3754
rect 191988 3726 192064 3754
rect 193184 3726 193260 3754
rect 194288 3726 194456 3754
rect 184952 480 184980 3726
rect 186148 480 186176 3726
rect 187344 480 187372 3726
rect 188540 480 188568 3726
rect 189736 480 189764 3726
rect 190840 480 190868 3726
rect 192036 480 192064 3726
rect 193232 480 193260 3726
rect 194428 480 194456 3726
rect 195440 3726 195512 3754
rect 196680 3754 196708 4012
rect 197784 3754 197812 4012
rect 198980 3754 199008 4012
rect 196680 3726 196848 3754
rect 197784 3726 197952 3754
rect 183714 190 183968 218
rect 183714 -960 183826 190
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195440 218 195468 3726
rect 196820 480 196848 3726
rect 197924 480 197952 3726
rect 198936 3726 199008 3754
rect 200084 3754 200112 4012
rect 201280 3754 201308 4012
rect 202476 3754 202504 4012
rect 203580 3754 203608 4012
rect 204776 3754 204804 4012
rect 205880 3754 205908 4012
rect 207076 3754 207104 4012
rect 208272 3754 208300 4012
rect 209376 3754 209404 4012
rect 210572 3754 210600 4012
rect 211676 3754 211704 4012
rect 212872 3754 212900 4012
rect 214068 3754 214096 4012
rect 215172 3754 215200 4012
rect 216368 3806 216396 4012
rect 216356 3800 216408 3806
rect 200084 3726 200344 3754
rect 201280 3726 201356 3754
rect 202476 3726 202736 3754
rect 203580 3726 203656 3754
rect 204776 3726 205128 3754
rect 205880 3726 206232 3754
rect 207076 3726 207152 3754
rect 208272 3726 208624 3754
rect 209376 3726 209728 3754
rect 210572 3726 211016 3754
rect 211676 3726 211752 3754
rect 212872 3726 213408 3754
rect 214068 3726 214512 3754
rect 215172 3726 215248 3754
rect 216356 3742 216408 3748
rect 216864 3800 216916 3806
rect 216864 3742 216916 3748
rect 217472 3754 217500 4012
rect 218668 3754 218696 4012
rect 219864 3754 219892 4012
rect 220968 3754 220996 4012
rect 222164 3806 222192 4012
rect 222152 3800 222204 3806
rect 195582 218 195694 480
rect 195440 190 195694 218
rect 195582 -960 195694 190
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198936 218 198964 3726
rect 200316 480 200344 3726
rect 199078 218 199190 480
rect 198936 190 199190 218
rect 199078 -960 199190 190
rect 200274 -960 200386 480
rect 201328 354 201356 3726
rect 202708 480 202736 3726
rect 201470 354 201582 480
rect 201328 326 201582 354
rect 201470 -960 201582 326
rect 202666 -960 202778 480
rect 203628 354 203656 3726
rect 205100 480 205128 3726
rect 206204 480 206232 3726
rect 203862 354 203974 480
rect 203628 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207124 354 207152 3726
rect 208596 480 208624 3726
rect 209700 626 209728 3726
rect 209700 598 209774 626
rect 209746 480 209774 598
rect 210988 480 211016 3726
rect 207358 354 207470 480
rect 207124 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209746 326 209862 480
rect 209750 -960 209862 326
rect 210946 -960 211058 480
rect 211724 354 211752 3726
rect 213380 480 213408 3726
rect 214484 480 214512 3726
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215220 354 215248 3726
rect 216876 480 216904 3742
rect 217472 3726 217640 3754
rect 218668 3726 219296 3754
rect 219864 3726 220032 3754
rect 220968 3726 221136 3754
rect 222152 3742 222204 3748
rect 222752 3800 222804 3806
rect 222752 3742 222804 3748
rect 223360 3754 223388 4012
rect 224464 3806 224492 4012
rect 224452 3800 224504 3806
rect 215638 354 215750 480
rect 215220 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 217612 354 217640 3726
rect 219268 480 219296 3726
rect 218030 354 218142 480
rect 217612 326 218142 354
rect 218030 -960 218142 326
rect 219226 -960 219338 480
rect 220004 354 220032 3726
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 3726
rect 222764 480 222792 3742
rect 223360 3726 223528 3754
rect 224452 3742 224504 3748
rect 225144 3800 225196 3806
rect 225144 3742 225196 3748
rect 225660 3754 225688 4012
rect 226764 3754 226792 4012
rect 227960 3754 227988 4012
rect 229156 3754 229184 4012
rect 230260 3806 230288 4012
rect 231456 3806 231484 4012
rect 232560 3806 232588 4012
rect 233756 3806 233784 4012
rect 230248 3800 230300 3806
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223500 354 223528 3726
rect 225156 480 225184 3742
rect 225660 3726 225920 3754
rect 226764 3726 227576 3754
rect 227960 3726 228312 3754
rect 229156 3726 229416 3754
rect 230248 3742 230300 3748
rect 231032 3800 231084 3806
rect 231032 3742 231084 3748
rect 231444 3800 231496 3806
rect 231444 3742 231496 3748
rect 232228 3800 232280 3806
rect 232228 3742 232280 3748
rect 232548 3800 232600 3806
rect 232548 3742 232600 3748
rect 233424 3800 233476 3806
rect 233424 3742 233476 3748
rect 233744 3800 233796 3806
rect 233744 3742 233796 3748
rect 234620 3800 234672 3806
rect 234620 3742 234672 3748
rect 234952 3754 234980 4012
rect 236056 3754 236084 4012
rect 237252 3806 237280 4012
rect 238356 3806 238384 4012
rect 239552 3806 239580 4012
rect 240748 3806 240776 4012
rect 241852 3806 241880 4012
rect 237240 3800 237292 3806
rect 223918 354 224030 480
rect 223500 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 225892 354 225920 3726
rect 227548 480 227576 3726
rect 226310 354 226422 480
rect 225892 326 226422 354
rect 226310 -960 226422 326
rect 227506 -960 227618 480
rect 228284 354 228312 3726
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 3726
rect 231044 480 231072 3742
rect 232240 480 232268 3742
rect 233436 480 233464 3742
rect 234632 480 234660 3742
rect 234952 3726 235856 3754
rect 236056 3726 236592 3754
rect 237240 3742 237292 3748
rect 238116 3800 238168 3806
rect 238116 3742 238168 3748
rect 238344 3800 238396 3806
rect 238344 3742 238396 3748
rect 239312 3800 239364 3806
rect 239312 3742 239364 3748
rect 239540 3800 239592 3806
rect 239540 3742 239592 3748
rect 240508 3800 240560 3806
rect 240508 3742 240560 3748
rect 240736 3800 240788 3806
rect 240736 3742 240788 3748
rect 241704 3800 241756 3806
rect 241704 3742 241756 3748
rect 241840 3800 241892 3806
rect 241840 3742 241892 3748
rect 242900 3800 242952 3806
rect 242900 3742 242952 3748
rect 243048 3754 243076 4012
rect 244152 3874 244180 4012
rect 244140 3868 244192 3874
rect 244140 3810 244192 3816
rect 245200 3868 245252 3874
rect 245200 3810 245252 3816
rect 235828 480 235856 3726
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 3726
rect 238128 480 238156 3742
rect 239324 480 239352 3742
rect 240520 480 240548 3742
rect 241716 480 241744 3742
rect 242912 480 242940 3742
rect 243048 3726 244136 3754
rect 244108 480 244136 3726
rect 245212 480 245240 3810
rect 245348 3806 245376 4012
rect 246544 3806 246572 4012
rect 247648 3942 247676 4012
rect 247636 3936 247688 3942
rect 247636 3878 247688 3884
rect 248604 3936 248656 3942
rect 248604 3878 248656 3884
rect 248844 3890 248872 4012
rect 245336 3800 245388 3806
rect 245336 3742 245388 3748
rect 246396 3800 246448 3806
rect 246396 3742 246448 3748
rect 246532 3800 246584 3806
rect 246532 3742 246584 3748
rect 247592 3800 247644 3806
rect 247592 3742 247644 3748
rect 246408 480 246436 3742
rect 247604 480 247632 3742
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 236982 -960 237094 326
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248616 354 248644 3878
rect 248844 3862 248920 3890
rect 248892 2854 248920 3862
rect 250040 3806 250068 4012
rect 251144 3890 251172 4012
rect 251100 3862 251172 3890
rect 250028 3800 250080 3806
rect 250028 3742 250080 3748
rect 251100 2854 251128 3862
rect 252340 3806 252368 4012
rect 253444 3890 253472 4012
rect 254640 3890 254668 4012
rect 253400 3862 253472 3890
rect 254596 3862 254668 3890
rect 251180 3800 251232 3806
rect 251180 3742 251232 3748
rect 252328 3800 252380 3806
rect 252328 3742 252380 3748
rect 248880 2848 248932 2854
rect 248880 2790 248932 2796
rect 249984 2848 250036 2854
rect 249984 2790 250036 2796
rect 251088 2848 251140 2854
rect 251088 2790 251140 2796
rect 249996 480 250024 2790
rect 251192 480 251220 3742
rect 253400 2922 253428 3862
rect 253480 3800 253532 3806
rect 253480 3742 253532 3748
rect 253388 2916 253440 2922
rect 253388 2858 253440 2864
rect 252376 2848 252428 2854
rect 252376 2790 252428 2796
rect 252388 480 252416 2790
rect 253492 480 253520 3742
rect 254596 2854 254624 3862
rect 255836 3806 255864 4012
rect 256940 3874 256968 4012
rect 256928 3868 256980 3874
rect 256928 3810 256980 3816
rect 258136 3806 258164 4012
rect 259240 3874 259268 4012
rect 258264 3868 258316 3874
rect 258264 3810 258316 3816
rect 259228 3868 259280 3874
rect 259228 3810 259280 3816
rect 255824 3800 255876 3806
rect 255824 3742 255876 3748
rect 257068 3800 257120 3806
rect 257068 3742 257120 3748
rect 258124 3800 258176 3806
rect 258124 3742 258176 3748
rect 254676 2916 254728 2922
rect 254676 2858 254728 2864
rect 254584 2848 254636 2854
rect 254584 2790 254636 2796
rect 254688 480 254716 2858
rect 255872 2848 255924 2854
rect 255872 2790 255924 2796
rect 255884 480 255912 2790
rect 257080 480 257108 3742
rect 258276 480 258304 3810
rect 260436 3806 260464 4012
rect 261632 3874 261660 4012
rect 260656 3868 260708 3874
rect 260656 3810 260708 3816
rect 261620 3868 261672 3874
rect 261620 3810 261672 3816
rect 259460 3800 259512 3806
rect 259460 3742 259512 3748
rect 260424 3800 260476 3806
rect 260424 3742 260476 3748
rect 259472 480 259500 3742
rect 260668 480 260696 3810
rect 262736 3806 262764 4012
rect 263932 3874 263960 4012
rect 262956 3868 263008 3874
rect 262956 3810 263008 3816
rect 263920 3868 263972 3874
rect 263920 3810 263972 3816
rect 261760 3800 261812 3806
rect 261760 3742 261812 3748
rect 262724 3800 262776 3806
rect 262724 3742 262776 3748
rect 261772 480 261800 3742
rect 262968 480 262996 3810
rect 265036 3806 265064 4012
rect 265348 3868 265400 3874
rect 265348 3810 265400 3816
rect 264152 3800 264204 3806
rect 264152 3742 264204 3748
rect 265024 3800 265076 3806
rect 265024 3742 265076 3748
rect 264164 480 264192 3742
rect 265360 480 265388 3810
rect 266232 3754 266260 4012
rect 267428 3806 267456 4012
rect 268532 3874 268560 4012
rect 268520 3868 268572 3874
rect 268520 3810 268572 3816
rect 269728 3806 269756 4012
rect 270832 3874 270860 4012
rect 270040 3868 270092 3874
rect 270040 3810 270092 3816
rect 270820 3868 270872 3874
rect 270820 3810 270872 3816
rect 266544 3800 266596 3806
rect 266232 3726 266308 3754
rect 266544 3742 266596 3748
rect 267416 3800 267468 3806
rect 267416 3742 267468 3748
rect 268844 3800 268896 3806
rect 268844 3742 268896 3748
rect 269716 3800 269768 3806
rect 269716 3742 269768 3748
rect 266280 1358 266308 3726
rect 266268 1352 266320 1358
rect 266268 1294 266320 1300
rect 266556 480 266584 3742
rect 267740 1352 267792 1358
rect 267740 1294 267792 1300
rect 267752 480 267780 1294
rect 268856 480 268884 3742
rect 270052 480 270080 3810
rect 272028 3806 272056 4012
rect 272432 3868 272484 3874
rect 272432 3810 272484 3816
rect 271236 3800 271288 3806
rect 271236 3742 271288 3748
rect 272016 3800 272068 3806
rect 272016 3742 272068 3748
rect 271248 480 271276 3742
rect 272444 480 272472 3810
rect 273224 3754 273252 4012
rect 273180 3726 273252 3754
rect 273628 3800 273680 3806
rect 273628 3742 273680 3748
rect 274328 3754 274356 4012
rect 275524 3874 275552 4012
rect 275512 3868 275564 3874
rect 275512 3810 275564 3816
rect 276720 3806 276748 4012
rect 277824 3874 277852 4012
rect 277124 3868 277176 3874
rect 277124 3810 277176 3816
rect 277812 3868 277864 3874
rect 277812 3810 277864 3816
rect 276708 3800 276760 3806
rect 273180 1358 273208 3726
rect 273168 1352 273220 1358
rect 273168 1294 273220 1300
rect 273640 480 273668 3742
rect 274328 3726 274404 3754
rect 276708 3742 276760 3748
rect 274376 746 274404 3726
rect 274824 1352 274876 1358
rect 274824 1294 274876 1300
rect 274364 740 274416 746
rect 274364 682 274416 688
rect 274836 480 274864 1294
rect 276020 740 276072 746
rect 276020 682 276072 688
rect 276032 480 276060 682
rect 277136 480 277164 3810
rect 279020 3806 279048 4012
rect 279516 3868 279568 3874
rect 279516 3810 279568 3816
rect 278320 3800 278372 3806
rect 278320 3742 278372 3748
rect 279008 3800 279060 3806
rect 279008 3742 279060 3748
rect 278332 480 278360 3742
rect 279528 480 279556 3810
rect 280124 3754 280152 4012
rect 280080 3726 280152 3754
rect 280712 3800 280764 3806
rect 280712 3742 280764 3748
rect 281320 3754 281348 4012
rect 282516 3754 282544 4012
rect 283620 3806 283648 4012
rect 284816 3874 284844 4012
rect 285920 3942 285948 4012
rect 285908 3936 285960 3942
rect 285908 3878 285960 3884
rect 284804 3868 284856 3874
rect 284804 3810 284856 3816
rect 286600 3868 286652 3874
rect 286600 3810 286652 3816
rect 283608 3800 283660 3806
rect 280080 1358 280108 3726
rect 280068 1352 280120 1358
rect 280068 1294 280120 1300
rect 280724 480 280752 3742
rect 281320 3726 281396 3754
rect 282516 3726 282592 3754
rect 283608 3742 283660 3748
rect 285404 3800 285456 3806
rect 285404 3742 285456 3748
rect 281368 1290 281396 3726
rect 282564 1358 282592 3726
rect 281908 1352 281960 1358
rect 281908 1294 281960 1300
rect 282552 1352 282604 1358
rect 282552 1294 282604 1300
rect 284300 1352 284352 1358
rect 284300 1294 284352 1300
rect 281356 1284 281408 1290
rect 281356 1226 281408 1232
rect 281920 480 281948 1294
rect 283104 1284 283156 1290
rect 283104 1226 283156 1232
rect 283116 480 283144 1226
rect 284312 480 284340 1294
rect 285416 480 285444 3742
rect 286612 480 286640 3810
rect 287116 3806 287144 4012
rect 287796 3936 287848 3942
rect 287796 3878 287848 3884
rect 287104 3800 287156 3806
rect 287104 3742 287156 3748
rect 287808 480 287836 3878
rect 288312 3754 288340 4012
rect 288992 3800 289044 3806
rect 288312 3726 288388 3754
rect 288992 3742 289044 3748
rect 289416 3754 289444 4012
rect 290612 3754 290640 4012
rect 291716 3806 291744 4012
rect 292912 3874 292940 4012
rect 292900 3868 292952 3874
rect 292900 3810 292952 3816
rect 294108 3806 294136 4012
rect 294880 3868 294932 3874
rect 294880 3810 294932 3816
rect 291704 3800 291756 3806
rect 288360 1358 288388 3726
rect 288348 1352 288400 1358
rect 288348 1294 288400 1300
rect 289004 480 289032 3742
rect 289416 3726 289492 3754
rect 290612 3726 290688 3754
rect 291704 3742 291756 3748
rect 293684 3800 293736 3806
rect 293684 3742 293736 3748
rect 294096 3800 294148 3806
rect 294096 3742 294148 3748
rect 289464 1290 289492 3726
rect 290188 1352 290240 1358
rect 290188 1294 290240 1300
rect 289452 1284 289504 1290
rect 289452 1226 289504 1232
rect 290200 480 290228 1294
rect 290660 610 290688 3726
rect 291384 1284 291436 1290
rect 291384 1226 291436 1232
rect 290648 604 290700 610
rect 290648 546 290700 552
rect 291396 480 291424 1226
rect 292580 604 292632 610
rect 292580 546 292632 552
rect 292592 480 292620 546
rect 293696 480 293724 3742
rect 294892 480 294920 3810
rect 295212 3754 295240 4012
rect 296076 3800 296128 3806
rect 295212 3726 295288 3754
rect 296076 3742 296128 3748
rect 296408 3754 296436 4012
rect 297512 3754 297540 4012
rect 298708 3806 298736 4012
rect 299904 3874 299932 4012
rect 299892 3868 299944 3874
rect 299892 3810 299944 3816
rect 301008 3806 301036 4012
rect 301964 3868 302016 3874
rect 301964 3810 302016 3816
rect 298696 3800 298748 3806
rect 295260 1358 295288 3726
rect 295248 1352 295300 1358
rect 295248 1294 295300 1300
rect 296088 480 296116 3742
rect 296408 3726 296484 3754
rect 297512 3726 297588 3754
rect 298696 3742 298748 3748
rect 300768 3800 300820 3806
rect 300768 3742 300820 3748
rect 300996 3800 301048 3806
rect 300996 3742 301048 3748
rect 296456 1290 296484 3726
rect 297560 1358 297588 3726
rect 297272 1352 297324 1358
rect 297272 1294 297324 1300
rect 297548 1352 297600 1358
rect 297548 1294 297600 1300
rect 299664 1352 299716 1358
rect 299664 1294 299716 1300
rect 296444 1284 296496 1290
rect 296444 1226 296496 1232
rect 297284 480 297312 1294
rect 298468 1284 298520 1290
rect 298468 1226 298520 1232
rect 298480 480 298508 1226
rect 299676 480 299704 1294
rect 300780 480 300808 3742
rect 301976 480 302004 3810
rect 302204 3754 302232 4012
rect 302160 3726 302232 3754
rect 303160 3800 303212 3806
rect 303160 3742 303212 3748
rect 303308 3754 303336 4012
rect 304504 3754 304532 4012
rect 305700 3754 305728 4012
rect 306804 3874 306832 4012
rect 306792 3868 306844 3874
rect 306792 3810 306844 3816
rect 308000 3806 308028 4012
rect 309048 3868 309100 3874
rect 309048 3810 309100 3816
rect 307988 3800 308040 3806
rect 302160 1358 302188 3726
rect 302148 1352 302200 1358
rect 302148 1294 302200 1300
rect 303172 480 303200 3742
rect 303308 3726 303384 3754
rect 304504 3726 304580 3754
rect 305700 3726 305776 3754
rect 307988 3742 308040 3748
rect 303356 1290 303384 3726
rect 304356 1352 304408 1358
rect 304356 1294 304408 1300
rect 303344 1284 303396 1290
rect 303344 1226 303396 1232
rect 304368 480 304396 1294
rect 304552 610 304580 3726
rect 305748 1358 305776 3726
rect 305736 1352 305788 1358
rect 305736 1294 305788 1300
rect 307944 1352 307996 1358
rect 307944 1294 307996 1300
rect 305552 1284 305604 1290
rect 305552 1226 305604 1232
rect 304540 604 304592 610
rect 304540 546 304592 552
rect 305564 480 305592 1226
rect 306748 604 306800 610
rect 306748 546 306800 552
rect 306760 480 306788 546
rect 307956 480 307984 1294
rect 309060 480 309088 3810
rect 309196 3754 309224 4012
rect 310300 3890 310328 4012
rect 311496 3890 311524 4012
rect 310300 3862 310376 3890
rect 311496 3862 311572 3890
rect 310244 3800 310296 3806
rect 309196 3726 309272 3754
rect 310244 3742 310296 3748
rect 309244 2854 309272 3726
rect 309232 2848 309284 2854
rect 309232 2790 309284 2796
rect 310256 480 310284 3742
rect 310348 1358 310376 3862
rect 311440 2848 311492 2854
rect 311440 2790 311492 2796
rect 310336 1352 310388 1358
rect 310336 1294 310388 1300
rect 311452 480 311480 2790
rect 311544 1222 311572 3862
rect 312600 3754 312628 4012
rect 312556 3726 312628 3754
rect 313796 3754 313824 4012
rect 314992 3754 315020 4012
rect 316096 3806 316124 4012
rect 316084 3800 316136 3806
rect 313796 3726 313872 3754
rect 314992 3726 315068 3754
rect 317292 3754 317320 4012
rect 316084 3742 316136 3748
rect 312556 1290 312584 3726
rect 313844 1358 313872 3726
rect 315040 2854 315068 3726
rect 317248 3726 317320 3754
rect 318396 3754 318424 4012
rect 318524 3800 318576 3806
rect 318396 3726 318472 3754
rect 318524 3742 318576 3748
rect 319592 3754 319620 4012
rect 320788 3754 320816 4012
rect 321892 3754 321920 4012
rect 323088 3806 323116 4012
rect 323076 3800 323128 3806
rect 315028 2848 315080 2854
rect 315028 2790 315080 2796
rect 317248 1358 317276 3726
rect 317328 2848 317380 2854
rect 317328 2790 317380 2796
rect 312636 1352 312688 1358
rect 312636 1294 312688 1300
rect 313832 1352 313884 1358
rect 313832 1294 313884 1300
rect 316224 1352 316276 1358
rect 316224 1294 316276 1300
rect 317236 1352 317288 1358
rect 317236 1294 317288 1300
rect 312544 1284 312596 1290
rect 312544 1226 312596 1232
rect 311532 1216 311584 1222
rect 311532 1158 311584 1164
rect 312648 480 312676 1294
rect 315028 1284 315080 1290
rect 315028 1226 315080 1232
rect 313832 1216 313884 1222
rect 313832 1158 313884 1164
rect 313844 480 313872 1158
rect 315040 480 315068 1226
rect 316236 480 316264 1294
rect 317340 480 317368 2790
rect 318444 1290 318472 3726
rect 318432 1284 318484 1290
rect 318432 1226 318484 1232
rect 318536 480 318564 3742
rect 319592 3726 319668 3754
rect 320788 3726 320864 3754
rect 321892 3726 321968 3754
rect 323076 3742 323128 3748
rect 324192 3754 324220 4012
rect 325388 3754 325416 4012
rect 325608 3800 325660 3806
rect 324192 3726 324268 3754
rect 325388 3726 325464 3754
rect 325608 3742 325660 3748
rect 326584 3754 326612 4012
rect 327688 3754 327716 4012
rect 328884 3754 328912 4012
rect 329988 3754 330016 4012
rect 331184 3754 331212 4012
rect 319640 1222 319668 3726
rect 319720 1352 319772 1358
rect 319720 1294 319772 1300
rect 319628 1216 319680 1222
rect 319628 1158 319680 1164
rect 319732 480 319760 1294
rect 320836 1154 320864 3726
rect 321940 1358 321968 3726
rect 321928 1352 321980 1358
rect 321928 1294 321980 1300
rect 324240 1290 324268 3726
rect 325436 1358 325464 3726
rect 324412 1352 324464 1358
rect 324412 1294 324464 1300
rect 325424 1352 325476 1358
rect 325424 1294 325476 1300
rect 320916 1284 320968 1290
rect 320916 1226 320968 1232
rect 324228 1284 324280 1290
rect 324228 1226 324280 1232
rect 320824 1148 320876 1154
rect 320824 1090 320876 1096
rect 320928 480 320956 1226
rect 322112 1216 322164 1222
rect 322112 1158 322164 1164
rect 322124 480 322152 1158
rect 323308 1148 323360 1154
rect 323308 1090 323360 1096
rect 323320 480 323348 1090
rect 324424 480 324452 1294
rect 325620 480 325648 3742
rect 326584 3726 326660 3754
rect 327688 3726 327764 3754
rect 328884 3726 328960 3754
rect 329988 3726 330064 3754
rect 326632 1222 326660 3726
rect 326804 1284 326856 1290
rect 326804 1226 326856 1232
rect 326620 1216 326672 1222
rect 326620 1158 326672 1164
rect 326816 480 326844 1226
rect 327736 1154 327764 3726
rect 328932 1358 328960 3726
rect 328000 1352 328052 1358
rect 328000 1294 328052 1300
rect 328920 1352 328972 1358
rect 328920 1294 328972 1300
rect 327724 1148 327776 1154
rect 327724 1090 327776 1096
rect 328012 480 328040 1294
rect 330036 1290 330064 3726
rect 331140 3726 331212 3754
rect 332380 3754 332408 4012
rect 333484 3754 333512 4012
rect 334680 3754 334708 4012
rect 335876 3754 335904 4012
rect 336980 3754 337008 4012
rect 338176 3754 338204 4012
rect 339280 3754 339308 4012
rect 340476 3754 340504 4012
rect 341672 3754 341700 4012
rect 342776 3754 342804 4012
rect 343972 3754 344000 4012
rect 345076 3754 345104 4012
rect 346272 3754 346300 4012
rect 347468 3754 347496 4012
rect 348572 3754 348600 4012
rect 349768 3754 349796 4012
rect 350872 3754 350900 4012
rect 352068 3754 352096 4012
rect 353264 3754 353292 4012
rect 332380 3726 332456 3754
rect 333484 3726 333560 3754
rect 334680 3726 334756 3754
rect 335876 3726 335952 3754
rect 336980 3726 337056 3754
rect 338176 3726 338252 3754
rect 339280 3726 339356 3754
rect 340476 3726 340552 3754
rect 341672 3726 341748 3754
rect 342776 3726 342852 3754
rect 343972 3726 344048 3754
rect 345076 3726 345152 3754
rect 346272 3726 346348 3754
rect 347468 3726 347544 3754
rect 348572 3726 348648 3754
rect 349768 3726 349844 3754
rect 350872 3726 350948 3754
rect 352068 3726 352144 3754
rect 330024 1284 330076 1290
rect 330024 1226 330076 1232
rect 331140 1222 331168 3726
rect 332428 1358 332456 3726
rect 331588 1352 331640 1358
rect 331588 1294 331640 1300
rect 332416 1352 332468 1358
rect 332416 1294 332468 1300
rect 329196 1216 329248 1222
rect 329196 1158 329248 1164
rect 331128 1216 331180 1222
rect 331128 1158 331180 1164
rect 329208 480 329236 1158
rect 330392 1148 330444 1154
rect 330392 1090 330444 1096
rect 330404 480 330432 1090
rect 331600 480 331628 1294
rect 332692 1284 332744 1290
rect 332692 1226 332744 1232
rect 332704 480 332732 1226
rect 333532 746 333560 3726
rect 334728 1290 334756 3726
rect 335924 1358 335952 3726
rect 335084 1352 335136 1358
rect 335084 1294 335136 1300
rect 335912 1352 335964 1358
rect 335912 1294 335964 1300
rect 334716 1284 334768 1290
rect 334716 1226 334768 1232
rect 333888 1216 333940 1222
rect 333888 1158 333940 1164
rect 333520 740 333572 746
rect 333520 682 333572 688
rect 333900 480 333928 1158
rect 335096 480 335124 1294
rect 337028 1222 337056 3726
rect 337476 1284 337528 1290
rect 337476 1226 337528 1232
rect 337016 1216 337068 1222
rect 337016 1158 337068 1164
rect 336280 740 336332 746
rect 336280 682 336332 688
rect 336292 480 336320 682
rect 337488 480 337516 1226
rect 338224 746 338252 3726
rect 339328 1358 339356 3726
rect 338672 1352 338724 1358
rect 338672 1294 338724 1300
rect 339316 1352 339368 1358
rect 339316 1294 339368 1300
rect 338212 740 338264 746
rect 338212 682 338264 688
rect 338684 480 338712 1294
rect 340524 1290 340552 3726
rect 340512 1284 340564 1290
rect 340512 1226 340564 1232
rect 341720 1222 341748 3726
rect 342168 1352 342220 1358
rect 342168 1294 342220 1300
rect 339868 1216 339920 1222
rect 339868 1158 339920 1164
rect 341708 1216 341760 1222
rect 341708 1158 341760 1164
rect 339880 480 339908 1158
rect 340972 740 341024 746
rect 340972 682 341024 688
rect 340984 480 341012 682
rect 342180 480 342208 1294
rect 342824 746 342852 3726
rect 344020 1290 344048 3726
rect 345124 1358 345152 3726
rect 345112 1352 345164 1358
rect 345112 1294 345164 1300
rect 343364 1284 343416 1290
rect 343364 1226 343416 1232
rect 344008 1284 344060 1290
rect 344008 1226 344060 1232
rect 342812 740 342864 746
rect 342812 682 342864 688
rect 343376 480 343404 1226
rect 344560 1216 344612 1222
rect 344560 1158 344612 1164
rect 344572 480 344600 1158
rect 346320 746 346348 3726
rect 346952 1284 347004 1290
rect 346952 1226 347004 1232
rect 345756 740 345808 746
rect 345756 682 345808 688
rect 346308 740 346360 746
rect 346308 682 346360 688
rect 345768 480 345796 682
rect 346964 480 346992 1226
rect 347516 882 347544 3726
rect 348056 1352 348108 1358
rect 348056 1294 348108 1300
rect 347504 876 347556 882
rect 347504 818 347556 824
rect 348068 480 348096 1294
rect 348620 1290 348648 3726
rect 349816 1358 349844 3726
rect 349804 1352 349856 1358
rect 349804 1294 349856 1300
rect 348608 1284 348660 1290
rect 348608 1226 348660 1232
rect 350448 876 350500 882
rect 350448 818 350500 824
rect 349252 740 349304 746
rect 349252 682 349304 688
rect 349264 480 349292 682
rect 350460 480 350488 818
rect 350920 746 350948 3726
rect 352116 1290 352144 3726
rect 353220 3726 353292 3754
rect 354368 3754 354396 4012
rect 355564 3754 355592 4012
rect 356668 3754 356696 4012
rect 357864 3754 357892 4012
rect 359060 3754 359088 4012
rect 360164 3754 360192 4012
rect 354368 3726 354444 3754
rect 355564 3726 355640 3754
rect 356668 3726 356744 3754
rect 357864 3726 357940 3754
rect 359060 3726 359136 3754
rect 353220 1358 353248 3726
rect 352840 1352 352892 1358
rect 352840 1294 352892 1300
rect 353208 1352 353260 1358
rect 353208 1294 353260 1300
rect 351644 1284 351696 1290
rect 351644 1226 351696 1232
rect 352104 1284 352156 1290
rect 352104 1226 352156 1232
rect 350908 740 350960 746
rect 350908 682 350960 688
rect 351656 480 351684 1226
rect 352852 480 352880 1294
rect 354036 740 354088 746
rect 354036 682 354088 688
rect 354048 480 354076 682
rect 248758 354 248870 480
rect 248616 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 354416 66 354444 3726
rect 355612 1290 355640 3726
rect 356716 1358 356744 3726
rect 356336 1352 356388 1358
rect 356336 1294 356388 1300
rect 356704 1352 356756 1358
rect 356704 1294 356756 1300
rect 355232 1284 355284 1290
rect 355232 1226 355284 1232
rect 355600 1284 355652 1290
rect 355600 1226 355652 1232
rect 355244 480 355272 1226
rect 356348 480 356376 1294
rect 357912 1222 357940 3726
rect 359108 1290 359136 3726
rect 360120 3726 360192 3754
rect 361360 3754 361388 4012
rect 362556 3754 362584 4012
rect 363660 3754 363688 4012
rect 364856 3754 364884 4012
rect 365960 3754 365988 4012
rect 367156 3754 367184 4012
rect 368352 3754 368380 4012
rect 369456 3754 369484 4012
rect 370652 3754 370680 4012
rect 371756 3754 371784 4012
rect 372952 3754 372980 4012
rect 374148 3754 374176 4012
rect 375252 3754 375280 4012
rect 376448 3754 376476 4012
rect 361360 3726 361436 3754
rect 362556 3726 362632 3754
rect 363660 3726 363736 3754
rect 364856 3726 364932 3754
rect 365960 3726 366036 3754
rect 367156 3726 367232 3754
rect 368352 3726 368428 3754
rect 369456 3726 369532 3754
rect 370652 3726 370728 3754
rect 371756 3726 371832 3754
rect 372952 3726 373028 3754
rect 374148 3726 374224 3754
rect 375252 3726 375328 3754
rect 359924 1352 359976 1358
rect 359924 1294 359976 1300
rect 358728 1284 358780 1290
rect 358728 1226 358780 1232
rect 359096 1284 359148 1290
rect 359096 1226 359148 1232
rect 357900 1216 357952 1222
rect 357900 1158 357952 1164
rect 358740 480 358768 1226
rect 359936 480 359964 1294
rect 360120 1154 360148 3726
rect 361120 1216 361172 1222
rect 361120 1158 361172 1164
rect 360108 1148 360160 1154
rect 360108 1090 360160 1096
rect 361132 480 361160 1158
rect 361408 882 361436 3726
rect 362604 1358 362632 3726
rect 362592 1352 362644 1358
rect 362592 1294 362644 1300
rect 363708 1290 363736 3726
rect 362316 1284 362368 1290
rect 362316 1226 362368 1232
rect 363696 1284 363748 1290
rect 363696 1226 363748 1232
rect 361396 876 361448 882
rect 361396 818 361448 824
rect 362328 480 362356 1226
rect 364904 1222 364932 3726
rect 365812 1352 365864 1358
rect 365812 1294 365864 1300
rect 364892 1216 364944 1222
rect 364892 1158 364944 1164
rect 363512 1148 363564 1154
rect 363512 1090 363564 1096
rect 363524 480 363552 1090
rect 364616 876 364668 882
rect 364616 818 364668 824
rect 364628 480 364656 818
rect 365824 480 365852 1294
rect 366008 746 366036 3726
rect 367204 1358 367232 3726
rect 367192 1352 367244 1358
rect 367192 1294 367244 1300
rect 367008 1284 367060 1290
rect 367008 1226 367060 1232
rect 365996 740 366048 746
rect 365996 682 366048 688
rect 367020 480 367048 1226
rect 368204 1216 368256 1222
rect 368204 1158 368256 1164
rect 368216 480 368244 1158
rect 368400 882 368428 3726
rect 368388 876 368440 882
rect 368388 818 368440 824
rect 369504 746 369532 3726
rect 370700 1358 370728 3726
rect 370596 1352 370648 1358
rect 370596 1294 370648 1300
rect 370688 1352 370740 1358
rect 370688 1294 370740 1300
rect 369400 740 369452 746
rect 369400 682 369452 688
rect 369492 740 369544 746
rect 369492 682 369544 688
rect 369412 480 369440 682
rect 370608 480 370636 1294
rect 371804 882 371832 3726
rect 373000 1290 373028 3726
rect 374092 1352 374144 1358
rect 374092 1294 374144 1300
rect 372988 1284 373040 1290
rect 372988 1226 373040 1232
rect 371700 876 371752 882
rect 371700 818 371752 824
rect 371792 876 371844 882
rect 371792 818 371844 824
rect 371712 480 371740 818
rect 372896 740 372948 746
rect 372896 682 372948 688
rect 372908 480 372936 682
rect 374104 480 374132 1294
rect 374196 1018 374224 3726
rect 375300 1222 375328 3726
rect 376404 3726 376476 3754
rect 377552 3754 377580 4012
rect 378748 3754 378776 4012
rect 379944 3754 379972 4012
rect 377552 3726 377628 3754
rect 378748 3726 378824 3754
rect 376404 1358 376432 3726
rect 376392 1352 376444 1358
rect 376392 1294 376444 1300
rect 377600 1290 377628 3726
rect 376484 1284 376536 1290
rect 376484 1226 376536 1232
rect 377588 1284 377640 1290
rect 377588 1226 377640 1232
rect 375288 1216 375340 1222
rect 375288 1158 375340 1164
rect 374184 1012 374236 1018
rect 374184 954 374236 960
rect 375288 876 375340 882
rect 375288 818 375340 824
rect 375300 480 375328 818
rect 376496 480 376524 1226
rect 378796 1086 378824 3726
rect 379900 3726 379972 3754
rect 381048 3754 381076 4012
rect 382244 3754 382272 4012
rect 381048 3726 381124 3754
rect 378876 1216 378928 1222
rect 378876 1158 378928 1164
rect 378784 1080 378836 1086
rect 378784 1022 378836 1028
rect 377680 1012 377732 1018
rect 377680 954 377732 960
rect 377692 480 377720 954
rect 378888 480 378916 1158
rect 379900 1018 379928 3726
rect 379980 1352 380032 1358
rect 379980 1294 380032 1300
rect 379888 1012 379940 1018
rect 379888 954 379940 960
rect 379992 480 380020 1294
rect 381096 1222 381124 3726
rect 382200 3726 382272 3754
rect 383348 3754 383376 4012
rect 384544 3754 384572 4012
rect 385740 3754 385768 4012
rect 386844 3754 386872 4012
rect 388040 3754 388068 4012
rect 389236 3754 389264 4012
rect 390340 3754 390368 4012
rect 391536 3754 391564 4012
rect 392640 3754 392668 4012
rect 393836 3754 393864 4012
rect 395032 3754 395060 4012
rect 396136 3754 396164 4012
rect 397332 3754 397360 4012
rect 398436 3754 398464 4012
rect 399632 3754 399660 4012
rect 400828 3754 400856 4012
rect 401932 3754 401960 4012
rect 403128 3754 403156 4012
rect 404232 3754 404260 4012
rect 405428 3754 405456 4012
rect 406624 3754 406652 4012
rect 407728 3754 407756 4012
rect 408924 3754 408952 4012
rect 410028 3754 410056 4012
rect 411224 3754 411252 4012
rect 383348 3726 383424 3754
rect 384544 3726 384620 3754
rect 385740 3726 385816 3754
rect 386844 3726 386920 3754
rect 388040 3726 388116 3754
rect 389236 3726 389312 3754
rect 390340 3726 390416 3754
rect 391536 3726 391612 3754
rect 392640 3726 392716 3754
rect 393836 3726 393912 3754
rect 395032 3726 395108 3754
rect 396136 3726 396212 3754
rect 397332 3726 397408 3754
rect 398436 3726 398512 3754
rect 399632 3726 399708 3754
rect 400828 3726 400904 3754
rect 401932 3726 402008 3754
rect 403128 3726 403204 3754
rect 404232 3726 404308 3754
rect 405428 3726 405504 3754
rect 406624 3726 406700 3754
rect 407728 3726 407804 3754
rect 408924 3726 409000 3754
rect 410028 3726 410104 3754
rect 381176 1284 381228 1290
rect 381176 1226 381228 1232
rect 381084 1216 381136 1222
rect 381084 1158 381136 1164
rect 381188 480 381216 1226
rect 382200 1154 382228 3726
rect 382188 1148 382240 1154
rect 382188 1090 382240 1096
rect 382372 1080 382424 1086
rect 382372 1022 382424 1028
rect 382384 480 382412 1022
rect 354404 60 354456 66
rect 354404 2 354456 8
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 82 357614 480
rect 357360 66 357614 82
rect 357348 60 357614 66
rect 357400 54 357614 60
rect 357348 2 357400 8
rect 357502 -960 357614 54
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383396 406 383424 3726
rect 383568 1012 383620 1018
rect 383568 954 383620 960
rect 383580 480 383608 954
rect 384592 882 384620 3726
rect 385788 1358 385816 3726
rect 385776 1352 385828 1358
rect 385776 1294 385828 1300
rect 384764 1216 384816 1222
rect 384764 1158 384816 1164
rect 384580 876 384632 882
rect 384580 818 384632 824
rect 384776 480 384804 1158
rect 385960 1148 386012 1154
rect 385960 1090 386012 1096
rect 385972 480 386000 1090
rect 386892 1086 386920 3726
rect 388088 1290 388116 3726
rect 388076 1284 388128 1290
rect 388076 1226 388128 1232
rect 389284 1154 389312 3726
rect 389456 1352 389508 1358
rect 389456 1294 389508 1300
rect 389272 1148 389324 1154
rect 389272 1090 389324 1096
rect 386880 1080 386932 1086
rect 386880 1022 386932 1028
rect 388260 876 388312 882
rect 388260 818 388312 824
rect 388272 480 388300 818
rect 389468 480 389496 1294
rect 390388 1222 390416 3726
rect 390376 1216 390428 1222
rect 390376 1158 390428 1164
rect 390652 1080 390704 1086
rect 390652 1022 390704 1028
rect 390664 480 390692 1022
rect 391584 882 391612 3726
rect 391848 1284 391900 1290
rect 391848 1226 391900 1232
rect 391572 876 391624 882
rect 391572 818 391624 824
rect 391860 480 391888 1226
rect 383384 400 383436 406
rect 383384 342 383436 348
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386788 400 386840 406
rect 387126 354 387238 480
rect 386840 348 387238 354
rect 386788 342 387238 348
rect 386800 326 387238 342
rect 387126 -960 387238 326
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392688 270 392716 3726
rect 393884 1290 393912 3726
rect 395080 1358 395108 3726
rect 395068 1352 395120 1358
rect 395068 1294 395120 1300
rect 393872 1284 393924 1290
rect 393872 1226 393924 1232
rect 394240 1216 394292 1222
rect 394240 1158 394292 1164
rect 393044 1148 393096 1154
rect 393044 1090 393096 1096
rect 393056 480 393084 1090
rect 394252 480 394280 1158
rect 396184 882 396212 3726
rect 397380 1154 397408 3726
rect 398484 1290 398512 3726
rect 399680 1358 399708 3726
rect 398932 1352 398984 1358
rect 398932 1294 398984 1300
rect 399668 1352 399720 1358
rect 399668 1294 399720 1300
rect 397736 1284 397788 1290
rect 397736 1226 397788 1232
rect 398472 1284 398524 1290
rect 398472 1226 398524 1232
rect 397368 1148 397420 1154
rect 397368 1090 397420 1096
rect 395344 876 395396 882
rect 395344 818 395396 824
rect 396172 876 396224 882
rect 396172 818 396224 824
rect 395356 480 395384 818
rect 397748 480 397776 1226
rect 398944 480 398972 1294
rect 400876 1222 400904 3726
rect 400864 1216 400916 1222
rect 400864 1158 400916 1164
rect 401324 1148 401376 1154
rect 401324 1090 401376 1096
rect 400128 876 400180 882
rect 400128 818 400180 824
rect 400140 480 400168 818
rect 401336 480 401364 1090
rect 392676 264 392728 270
rect 392676 206 392728 212
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396172 264 396224 270
rect 396510 218 396622 480
rect 396224 212 396622 218
rect 396172 206 396622 212
rect 396184 190 396622 206
rect 396510 -960 396622 190
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 401980 66 402008 3726
rect 403176 1290 403204 3726
rect 403624 1352 403676 1358
rect 403624 1294 403676 1300
rect 402520 1284 402572 1290
rect 402520 1226 402572 1232
rect 403164 1284 403216 1290
rect 403164 1226 403216 1232
rect 402532 480 402560 1226
rect 403636 480 403664 1294
rect 404280 1154 404308 3726
rect 405476 1358 405504 3726
rect 405464 1352 405516 1358
rect 405464 1294 405516 1300
rect 404820 1216 404872 1222
rect 404820 1158 404872 1164
rect 404268 1148 404320 1154
rect 404268 1090 404320 1096
rect 404832 480 404860 1158
rect 406672 882 406700 3726
rect 407212 1284 407264 1290
rect 407212 1226 407264 1232
rect 406660 876 406712 882
rect 406660 818 406712 824
rect 407224 480 407252 1226
rect 407776 1222 407804 3726
rect 407764 1216 407816 1222
rect 407764 1158 407816 1164
rect 408972 1154 409000 3726
rect 409604 1352 409656 1358
rect 409604 1294 409656 1300
rect 408408 1148 408460 1154
rect 408408 1090 408460 1096
rect 408960 1148 409012 1154
rect 408960 1090 409012 1096
rect 408420 480 408448 1090
rect 409616 480 409644 1294
rect 410076 1290 410104 3726
rect 411180 3726 411252 3754
rect 412420 3754 412448 4012
rect 413524 3754 413552 4012
rect 414720 3754 414748 4012
rect 415916 3754 415944 4012
rect 417020 3754 417048 4012
rect 418216 3754 418244 4012
rect 419320 3754 419348 4012
rect 420516 3754 420544 4012
rect 421712 3754 421740 4012
rect 422816 3754 422844 4012
rect 424012 3754 424040 4012
rect 425116 3754 425144 4012
rect 426312 3754 426340 4012
rect 427508 3754 427536 4012
rect 428612 3754 428640 4012
rect 429808 3754 429836 4012
rect 430912 3754 430940 4012
rect 432108 3754 432136 4012
rect 433304 3754 433332 4012
rect 434408 3754 434436 4012
rect 412420 3726 412496 3754
rect 413524 3726 413600 3754
rect 414720 3726 414796 3754
rect 415916 3726 415992 3754
rect 417020 3726 417096 3754
rect 418216 3726 418292 3754
rect 419320 3726 419396 3754
rect 420516 3726 420592 3754
rect 421712 3726 421788 3754
rect 422816 3726 422892 3754
rect 424012 3726 424088 3754
rect 425116 3726 425192 3754
rect 426312 3726 426388 3754
rect 427508 3726 427584 3754
rect 428612 3726 428688 3754
rect 429808 3726 429884 3754
rect 430912 3726 431080 3754
rect 432108 3726 432184 3754
rect 411180 2854 411208 3726
rect 411168 2848 411220 2854
rect 411168 2790 411220 2796
rect 410064 1284 410116 1290
rect 410064 1226 410116 1232
rect 411904 1216 411956 1222
rect 411904 1158 411956 1164
rect 410800 876 410852 882
rect 410800 818 410852 824
rect 410812 480 410840 818
rect 411916 480 411944 1158
rect 401968 60 402020 66
rect 401968 2 402020 8
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 82 406098 480
rect 405986 66 406240 82
rect 405986 60 406252 66
rect 405986 54 406200 60
rect 405986 -960 406098 54
rect 406200 2 406252 8
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412468 270 412496 3726
rect 413572 1222 413600 3726
rect 414296 1284 414348 1290
rect 414296 1226 414348 1232
rect 413560 1216 413612 1222
rect 413560 1158 413612 1164
rect 413100 1148 413152 1154
rect 413100 1090 413152 1096
rect 413112 480 413140 1090
rect 414308 480 414336 1226
rect 414768 1018 414796 3726
rect 415492 2848 415544 2854
rect 415492 2790 415544 2796
rect 414756 1012 414808 1018
rect 414756 954 414808 960
rect 415504 480 415532 2790
rect 415964 1358 415992 3726
rect 415952 1352 416004 1358
rect 415952 1294 416004 1300
rect 417068 882 417096 3726
rect 418264 1290 418292 3726
rect 418252 1284 418304 1290
rect 418252 1226 418304 1232
rect 419368 1222 419396 3726
rect 420184 1352 420236 1358
rect 420184 1294 420236 1300
rect 417884 1216 417936 1222
rect 417884 1158 417936 1164
rect 419356 1216 419408 1222
rect 419356 1158 419408 1164
rect 417056 876 417108 882
rect 417056 818 417108 824
rect 417896 480 417924 1158
rect 418988 1012 419040 1018
rect 418988 954 419040 960
rect 419000 480 419028 954
rect 420196 480 420224 1294
rect 420564 1154 420592 3726
rect 420552 1148 420604 1154
rect 420552 1090 420604 1096
rect 421380 876 421432 882
rect 421380 818 421432 824
rect 421392 480 421420 818
rect 412456 264 412508 270
rect 412456 206 412508 212
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 218 416770 480
rect 416872 264 416924 270
rect 416658 212 416872 218
rect 416658 206 416924 212
rect 416658 190 416912 206
rect 416658 -960 416770 190
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 421760 270 421788 3726
rect 422576 1284 422628 1290
rect 422576 1226 422628 1232
rect 422588 480 422616 1226
rect 422864 1018 422892 3726
rect 424060 1290 424088 3726
rect 424048 1284 424100 1290
rect 424048 1226 424100 1232
rect 423404 1216 423456 1222
rect 423404 1158 423456 1164
rect 422852 1012 422904 1018
rect 422852 954 422904 960
rect 421748 264 421800 270
rect 421748 206 421800 212
rect 422546 -960 422658 480
rect 423416 354 423444 1158
rect 424968 1148 425020 1154
rect 424968 1090 425020 1096
rect 424980 480 425008 1090
rect 425164 1086 425192 3726
rect 426360 1222 426388 3726
rect 427556 1358 427584 3726
rect 427544 1352 427596 1358
rect 427544 1294 427596 1300
rect 428464 1284 428516 1290
rect 428464 1226 428516 1232
rect 426348 1216 426400 1222
rect 426348 1158 426400 1164
rect 425152 1080 425204 1086
rect 425152 1022 425204 1028
rect 427268 1012 427320 1018
rect 427268 954 427320 960
rect 427280 480 427308 954
rect 428476 480 428504 1226
rect 428660 1154 428688 3726
rect 428648 1148 428700 1154
rect 428648 1090 428700 1096
rect 429660 1080 429712 1086
rect 429660 1022 429712 1028
rect 429672 480 429700 1022
rect 429856 882 429884 3726
rect 430856 1216 430908 1222
rect 430856 1158 430908 1164
rect 429844 876 429896 882
rect 429844 818 429896 824
rect 430868 480 430896 1158
rect 423742 354 423854 480
rect 423416 326 423854 354
rect 423742 -960 423854 326
rect 424938 -960 425050 480
rect 425796 264 425848 270
rect 426134 218 426246 480
rect 425848 212 426246 218
rect 425796 206 426246 212
rect 425808 190 426246 206
rect 426134 -960 426246 190
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 431052 134 431080 3726
rect 431868 1352 431920 1358
rect 431868 1294 431920 1300
rect 431880 354 431908 1294
rect 432156 1018 432184 3726
rect 433260 3726 433332 3754
rect 434364 3726 434436 3754
rect 435604 3754 435632 4012
rect 436708 3754 436736 4012
rect 437904 3754 437932 4012
rect 439100 3754 439128 4012
rect 440204 3754 440232 4012
rect 435604 3726 435680 3754
rect 436708 3726 436784 3754
rect 437904 3726 437980 3754
rect 439100 3726 439176 3754
rect 433260 1358 433288 3726
rect 433248 1352 433300 1358
rect 433248 1294 433300 1300
rect 433248 1148 433300 1154
rect 433248 1090 433300 1096
rect 432144 1012 432196 1018
rect 432144 954 432196 960
rect 433260 480 433288 1090
rect 434364 814 434392 3726
rect 435652 1290 435680 3726
rect 435640 1284 435692 1290
rect 435640 1226 435692 1232
rect 436756 1154 436784 3726
rect 437848 1352 437900 1358
rect 437848 1294 437900 1300
rect 436744 1148 436796 1154
rect 436744 1090 436796 1096
rect 436744 1012 436796 1018
rect 436744 954 436796 960
rect 434444 876 434496 882
rect 434444 818 434496 824
rect 434352 808 434404 814
rect 434352 750 434404 756
rect 434456 480 434484 818
rect 436756 480 436784 954
rect 437860 762 437888 1294
rect 437952 950 437980 3726
rect 439148 1086 439176 3726
rect 440160 3726 440232 3754
rect 441400 3754 441428 4012
rect 442596 3754 442624 4012
rect 443700 3754 443728 4012
rect 444896 3754 444924 4012
rect 446000 3754 446028 4012
rect 447196 3754 447224 4012
rect 448392 3754 448420 4012
rect 449496 3754 449524 4012
rect 450692 3754 450720 4012
rect 451796 3754 451824 4012
rect 452992 3754 453020 4012
rect 454188 3754 454216 4012
rect 455292 3754 455320 4012
rect 456488 3754 456516 4012
rect 457592 3754 457620 4012
rect 458788 3754 458816 4012
rect 459984 3754 460012 4012
rect 461088 3754 461116 4012
rect 462284 3754 462312 4012
rect 441400 3726 441476 3754
rect 442596 3726 442672 3754
rect 443700 3726 443776 3754
rect 444896 3726 444972 3754
rect 446000 3726 446076 3754
rect 447196 3726 447272 3754
rect 448392 3726 448468 3754
rect 449496 3726 449572 3754
rect 450692 3726 450768 3754
rect 451796 3726 451872 3754
rect 452992 3726 453068 3754
rect 454188 3726 454264 3754
rect 455292 3726 455368 3754
rect 456488 3726 456564 3754
rect 457592 3726 457668 3754
rect 458788 3726 458864 3754
rect 459984 3726 460060 3754
rect 461088 3726 461164 3754
rect 440160 2854 440188 3726
rect 440148 2848 440200 2854
rect 440148 2790 440200 2796
rect 439964 1284 440016 1290
rect 439964 1226 440016 1232
rect 439136 1080 439188 1086
rect 439136 1022 439188 1028
rect 437940 944 437992 950
rect 437940 886 437992 892
rect 439136 808 439188 814
rect 437860 734 437980 762
rect 439136 750 439188 756
rect 437952 480 437980 734
rect 439148 480 439176 750
rect 432022 354 432134 480
rect 431880 326 432134 354
rect 431040 128 431092 134
rect 431040 70 431092 76
rect 432022 -960 432134 326
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435180 128 435232 134
rect 435518 82 435630 480
rect 435232 76 435630 82
rect 435180 70 435630 76
rect 435192 54 435630 70
rect 435518 -960 435630 54
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 439976 354 440004 1226
rect 441448 1222 441476 3726
rect 442644 1358 442672 3726
rect 442632 1352 442684 1358
rect 442632 1294 442684 1300
rect 441436 1216 441488 1222
rect 441436 1158 441488 1164
rect 441528 1148 441580 1154
rect 441528 1090 441580 1096
rect 441540 480 441568 1090
rect 442632 944 442684 950
rect 442632 886 442684 892
rect 442644 480 442672 886
rect 443748 882 443776 3726
rect 444944 1290 444972 3726
rect 445024 2848 445076 2854
rect 445024 2790 445076 2796
rect 444932 1284 444984 1290
rect 444932 1226 444984 1232
rect 443828 1080 443880 1086
rect 443828 1022 443880 1028
rect 443736 876 443788 882
rect 443736 818 443788 824
rect 443840 480 443868 1022
rect 445036 480 445064 2790
rect 446048 1222 446076 3726
rect 445852 1216 445904 1222
rect 445852 1158 445904 1164
rect 446036 1216 446088 1222
rect 446036 1158 446088 1164
rect 440302 354 440414 480
rect 439976 326 440414 354
rect 440302 -960 440414 326
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445864 354 445892 1158
rect 447244 1086 447272 3726
rect 448440 1358 448468 3726
rect 449544 2854 449572 3726
rect 449532 2848 449584 2854
rect 449532 2790 449584 2796
rect 447416 1352 447468 1358
rect 447416 1294 447468 1300
rect 448428 1352 448480 1358
rect 448428 1294 448480 1300
rect 447232 1080 447284 1086
rect 447232 1022 447284 1028
rect 447428 480 447456 1294
rect 450740 1290 450768 3726
rect 449808 1284 449860 1290
rect 449808 1226 449860 1232
rect 450728 1284 450780 1290
rect 450728 1226 450780 1232
rect 448244 876 448296 882
rect 448244 818 448296 824
rect 446190 354 446302 480
rect 445864 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448256 354 448284 818
rect 449820 480 449848 1226
rect 450912 1216 450964 1222
rect 450912 1158 450964 1164
rect 450924 480 450952 1158
rect 451844 882 451872 3726
rect 452108 1080 452160 1086
rect 452108 1022 452160 1028
rect 451832 876 451884 882
rect 451832 818 451884 824
rect 452120 480 452148 1022
rect 453040 1018 453068 3726
rect 453304 1352 453356 1358
rect 453304 1294 453356 1300
rect 453028 1012 453080 1018
rect 453028 954 453080 960
rect 453316 480 453344 1294
rect 454236 1154 454264 3726
rect 454500 2848 454552 2854
rect 454500 2790 454552 2796
rect 454224 1148 454276 1154
rect 454224 1090 454276 1096
rect 454512 480 454540 2790
rect 455340 1086 455368 3726
rect 456536 1290 456564 3726
rect 455696 1284 455748 1290
rect 455696 1226 455748 1232
rect 456524 1284 456576 1290
rect 456524 1226 456576 1232
rect 455328 1080 455380 1086
rect 455328 1022 455380 1028
rect 455708 480 455736 1226
rect 457640 1222 457668 3726
rect 458836 1358 458864 3726
rect 458824 1352 458876 1358
rect 458824 1294 458876 1300
rect 457628 1216 457680 1222
rect 457628 1158 457680 1164
rect 459192 1148 459244 1154
rect 459192 1090 459244 1096
rect 458088 1012 458140 1018
rect 458088 954 458140 960
rect 456524 876 456576 882
rect 456524 818 456576 824
rect 448582 354 448694 480
rect 448256 326 448694 354
rect 448582 -960 448694 326
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456536 354 456564 818
rect 458100 480 458128 954
rect 459204 480 459232 1090
rect 456862 354 456974 480
rect 456536 326 456974 354
rect 456862 -960 456974 326
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460032 134 460060 3726
rect 461136 1154 461164 3726
rect 462240 3726 462312 3754
rect 463388 3754 463416 4012
rect 464584 3754 464612 4012
rect 465780 3754 465808 4012
rect 466884 3754 466912 4012
rect 468080 3754 468108 4012
rect 469276 3754 469304 4012
rect 470380 3754 470408 4012
rect 471576 3754 471604 4012
rect 472680 3754 472708 4012
rect 473876 3754 473904 4012
rect 475072 3754 475100 4012
rect 476176 3754 476204 4012
rect 477372 3754 477400 4012
rect 478476 3754 478504 4012
rect 479672 3754 479700 4012
rect 480868 3754 480896 4012
rect 481972 3754 482000 4012
rect 483168 3754 483196 4012
rect 484272 3754 484300 4012
rect 485468 3754 485496 4012
rect 486664 3754 486692 4012
rect 487768 3754 487796 4012
rect 488964 3754 488992 4012
rect 490068 3754 490096 4012
rect 491264 3754 491292 4012
rect 463388 3726 463464 3754
rect 464584 3726 464660 3754
rect 465780 3726 465856 3754
rect 466884 3726 466960 3754
rect 468080 3726 468156 3754
rect 469276 3726 469352 3754
rect 470380 3726 470456 3754
rect 471576 3726 471652 3754
rect 472680 3726 472756 3754
rect 473876 3726 473952 3754
rect 475072 3726 475148 3754
rect 476176 3726 476252 3754
rect 477372 3726 477448 3754
rect 478476 3726 478552 3754
rect 479672 3726 479748 3754
rect 480868 3726 480944 3754
rect 481972 3726 482048 3754
rect 483168 3726 483244 3754
rect 484272 3726 484348 3754
rect 485468 3726 485544 3754
rect 486664 3726 486740 3754
rect 487768 3726 487844 3754
rect 488964 3726 489040 3754
rect 490068 3726 490144 3754
rect 462240 1290 462268 3726
rect 461584 1284 461636 1290
rect 461584 1226 461636 1232
rect 462228 1284 462280 1290
rect 462228 1226 462280 1232
rect 461124 1148 461176 1154
rect 461124 1090 461176 1096
rect 460112 1080 460164 1086
rect 460112 1022 460164 1028
rect 460124 354 460152 1022
rect 461596 480 461624 1226
rect 462412 1216 462464 1222
rect 462412 1158 462464 1164
rect 460358 354 460470 480
rect 460124 326 460470 354
rect 460020 128 460072 134
rect 460020 70 460072 76
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462424 354 462452 1158
rect 463436 882 463464 3726
rect 463976 1352 464028 1358
rect 463976 1294 464028 1300
rect 463424 876 463476 882
rect 463424 818 463476 824
rect 463988 480 464016 1294
rect 464632 1018 464660 3726
rect 465828 1222 465856 3726
rect 465816 1216 465868 1222
rect 465816 1158 465868 1164
rect 466276 1148 466328 1154
rect 466276 1090 466328 1096
rect 464620 1012 464672 1018
rect 464620 954 464672 960
rect 466288 480 466316 1090
rect 466932 1086 466960 3726
rect 468128 1358 468156 3726
rect 468116 1352 468168 1358
rect 468116 1294 468168 1300
rect 467472 1284 467524 1290
rect 467472 1226 467524 1232
rect 466920 1080 466972 1086
rect 466920 1022 466972 1028
rect 467484 480 467512 1226
rect 468668 876 468720 882
rect 468668 818 468720 824
rect 468680 480 468708 818
rect 462750 354 462862 480
rect 462424 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 464988 128 465040 134
rect 465142 82 465254 480
rect 465040 76 465254 82
rect 464988 70 465254 76
rect 465000 54 465254 70
rect 465142 -960 465254 54
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469324 270 469352 3726
rect 469864 1012 469916 1018
rect 469864 954 469916 960
rect 469876 480 469904 954
rect 469312 264 469364 270
rect 469312 206 469364 212
rect 469834 -960 469946 480
rect 470428 134 470456 3726
rect 471624 1290 471652 3726
rect 471612 1284 471664 1290
rect 471612 1226 471664 1232
rect 470692 1216 470744 1222
rect 470692 1158 470744 1164
rect 470704 354 470732 1158
rect 472728 1154 472756 3726
rect 473084 1352 473136 1358
rect 473084 1294 473136 1300
rect 472716 1148 472768 1154
rect 472716 1090 472768 1096
rect 472256 1080 472308 1086
rect 472256 1022 472308 1028
rect 472268 480 472296 1022
rect 471030 354 471142 480
rect 470704 326 471142 354
rect 470416 128 470468 134
rect 470416 70 470468 76
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473096 354 473124 1294
rect 473924 1018 473952 3726
rect 475120 1222 475148 3726
rect 475108 1216 475160 1222
rect 475108 1158 475160 1164
rect 473912 1012 473964 1018
rect 473912 954 473964 960
rect 476224 882 476252 3726
rect 476580 1284 476632 1290
rect 476580 1226 476632 1232
rect 476212 876 476264 882
rect 476212 818 476264 824
rect 473422 354 473534 480
rect 473096 326 473534 354
rect 473422 -960 473534 326
rect 474188 264 474240 270
rect 474526 218 474638 480
rect 474240 212 474638 218
rect 474188 206 474638 212
rect 474200 190 474638 206
rect 474526 -960 474638 190
rect 475722 82 475834 480
rect 476592 354 476620 1226
rect 477420 1086 477448 3726
rect 478524 2854 478552 3726
rect 478512 2848 478564 2854
rect 478512 2790 478564 2796
rect 479720 1290 479748 3726
rect 480916 1358 480944 3726
rect 480904 1352 480956 1358
rect 480904 1294 480956 1300
rect 479708 1284 479760 1290
rect 479708 1226 479760 1232
rect 482020 1222 482048 3726
rect 480536 1216 480588 1222
rect 480536 1158 480588 1164
rect 482008 1216 482060 1222
rect 482008 1158 482060 1164
rect 478144 1148 478196 1154
rect 478144 1090 478196 1096
rect 477408 1080 477460 1086
rect 477408 1022 477460 1028
rect 478156 480 478184 1090
rect 479340 1012 479392 1018
rect 479340 954 479392 960
rect 479352 480 479380 954
rect 480548 480 480576 1158
rect 482468 1080 482520 1086
rect 482468 1022 482520 1028
rect 481364 876 481416 882
rect 481364 818 481416 824
rect 476918 354 477030 480
rect 476592 326 477030 354
rect 475936 128 475988 134
rect 475722 76 475936 82
rect 475722 70 475988 76
rect 475722 54 475976 70
rect 475722 -960 475834 54
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481376 354 481404 818
rect 481702 354 481814 480
rect 481376 326 481814 354
rect 482480 354 482508 1022
rect 483216 950 483244 3726
rect 484032 2848 484084 2854
rect 484032 2790 484084 2796
rect 483204 944 483256 950
rect 483204 886 483256 892
rect 484044 480 484072 2790
rect 484320 1018 484348 3726
rect 484860 1284 484912 1290
rect 484860 1226 484912 1232
rect 484308 1012 484360 1018
rect 484308 954 484360 960
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 481702 -960 481814 326
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484872 354 484900 1226
rect 485516 1086 485544 3726
rect 486424 1352 486476 1358
rect 486424 1294 486476 1300
rect 485504 1080 485556 1086
rect 485504 1022 485556 1028
rect 486436 480 486464 1294
rect 486712 1154 486740 3726
rect 487816 1358 487844 3726
rect 487804 1352 487856 1358
rect 487804 1294 487856 1300
rect 489012 1290 489040 3726
rect 489000 1284 489052 1290
rect 489000 1226 489052 1232
rect 487252 1216 487304 1222
rect 487252 1158 487304 1164
rect 486700 1148 486752 1154
rect 486700 1090 486752 1096
rect 485198 354 485310 480
rect 484872 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487264 354 487292 1158
rect 490116 1018 490144 3726
rect 491220 3726 491292 3754
rect 492460 3754 492488 4012
rect 493564 3754 493592 4012
rect 494760 3754 494788 4012
rect 495956 3754 495984 4012
rect 497060 3754 497088 4012
rect 498256 3754 498284 4012
rect 499360 3754 499388 4012
rect 500556 3754 500584 4012
rect 501752 3754 501780 4012
rect 492460 3726 492536 3754
rect 493564 3726 493640 3754
rect 494760 3726 494836 3754
rect 495956 3726 496032 3754
rect 497060 3726 497136 3754
rect 498256 3726 498332 3754
rect 490748 1080 490800 1086
rect 490748 1022 490800 1028
rect 489920 1012 489972 1018
rect 489920 954 489972 960
rect 490104 1012 490156 1018
rect 490104 954 490156 960
rect 488816 944 488868 950
rect 488816 886 488868 892
rect 488828 480 488856 886
rect 489932 480 489960 954
rect 487590 354 487702 480
rect 487264 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 1022
rect 491220 950 491248 3726
rect 492508 1222 492536 3726
rect 493140 1352 493192 1358
rect 493140 1294 493192 1300
rect 492496 1216 492548 1222
rect 492496 1158 492548 1164
rect 492312 1148 492364 1154
rect 492312 1090 492364 1096
rect 491208 944 491260 950
rect 491208 886 491260 892
rect 492324 480 492352 1090
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493152 354 493180 1294
rect 493612 1154 493640 3726
rect 494704 1284 494756 1290
rect 494704 1226 494756 1232
rect 493600 1148 493652 1154
rect 493600 1090 493652 1096
rect 494716 480 494744 1226
rect 494808 1086 494836 3726
rect 494796 1080 494848 1086
rect 494796 1022 494848 1028
rect 496004 1018 496032 3726
rect 497108 1358 497136 3726
rect 497096 1352 497148 1358
rect 497096 1294 497148 1300
rect 498304 1290 498332 3726
rect 499224 3726 499388 3754
rect 500512 3726 500584 3754
rect 501708 3726 501780 3754
rect 502856 3754 502884 4012
rect 504052 3754 504080 4012
rect 505156 3754 505184 4012
rect 506352 3754 506380 4012
rect 507548 3754 507576 4012
rect 502856 3726 502932 3754
rect 504052 3726 504128 3754
rect 505156 3726 505232 3754
rect 498292 1284 498344 1290
rect 498292 1226 498344 1232
rect 498200 1216 498252 1222
rect 498200 1158 498252 1164
rect 495532 1012 495584 1018
rect 495532 954 495584 960
rect 495992 1012 496044 1018
rect 495992 954 496044 960
rect 493478 354 493590 480
rect 493152 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495544 354 495572 954
rect 497096 944 497148 950
rect 497096 886 497148 892
rect 497108 480 497136 886
rect 498212 480 498240 1158
rect 495870 354 495982 480
rect 495544 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499224 66 499252 3726
rect 500512 1154 500540 3726
rect 499396 1148 499448 1154
rect 499396 1090 499448 1096
rect 500500 1148 500552 1154
rect 500500 1090 500552 1096
rect 499408 480 499436 1090
rect 501708 1086 501736 3726
rect 500592 1080 500644 1086
rect 500592 1022 500644 1028
rect 501696 1080 501748 1086
rect 501696 1022 501748 1028
rect 500604 480 500632 1022
rect 502904 1018 502932 3726
rect 504100 1358 504128 3726
rect 502984 1352 503036 1358
rect 502984 1294 503036 1300
rect 504088 1352 504140 1358
rect 504088 1294 504140 1300
rect 501788 1012 501840 1018
rect 501788 954 501840 960
rect 502892 1012 502944 1018
rect 502892 954 502944 960
rect 501800 480 501828 954
rect 502996 480 503024 1294
rect 503812 1284 503864 1290
rect 503812 1226 503864 1232
rect 499212 60 499264 66
rect 499212 2 499264 8
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503824 354 503852 1226
rect 505204 1222 505232 3726
rect 506308 3726 506380 3754
rect 507504 3726 507576 3754
rect 508652 3754 508680 4012
rect 509848 3754 509876 4012
rect 510952 3754 510980 4012
rect 512148 3754 512176 4012
rect 513344 3754 513372 4012
rect 508652 3726 508728 3754
rect 509848 3726 509924 3754
rect 510952 3726 511028 3754
rect 512148 3726 512224 3754
rect 505192 1216 505244 1222
rect 505192 1158 505244 1164
rect 504150 354 504262 480
rect 503824 326 504262 354
rect 504150 -960 504262 326
rect 505346 82 505458 480
rect 505346 66 505600 82
rect 506308 66 506336 3726
rect 506480 1148 506532 1154
rect 506480 1090 506532 1096
rect 506492 480 506520 1090
rect 507308 1080 507360 1086
rect 507308 1022 507360 1028
rect 505346 60 505612 66
rect 505346 54 505560 60
rect 505346 -960 505458 54
rect 505560 2 505612 8
rect 506296 60 506348 66
rect 506296 2 506348 8
rect 506450 -960 506562 480
rect 507320 354 507348 1022
rect 507504 474 507532 3726
rect 507492 468 507544 474
rect 507492 410 507544 416
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 508700 270 508728 3726
rect 509896 1358 509924 3726
rect 509700 1352 509752 1358
rect 509700 1294 509752 1300
rect 509884 1352 509936 1358
rect 509884 1294 509936 1300
rect 508872 1012 508924 1018
rect 508872 954 508924 960
rect 508884 480 508912 954
rect 508688 264 508740 270
rect 508688 206 508740 212
rect 508842 -960 508954 480
rect 509712 354 509740 1294
rect 511000 1290 511028 3726
rect 510988 1284 511040 1290
rect 510988 1226 511040 1232
rect 511264 1216 511316 1222
rect 511264 1158 511316 1164
rect 511276 480 511304 1158
rect 512196 1154 512224 3726
rect 513300 3726 513372 3754
rect 514448 3754 514476 4012
rect 515644 3754 515672 4012
rect 516748 3754 516776 4012
rect 517944 3754 517972 4012
rect 519140 3754 519168 4012
rect 520244 3754 520272 4012
rect 514448 3726 514524 3754
rect 515644 3726 515720 3754
rect 516748 3726 516824 3754
rect 517944 3726 518020 3754
rect 519140 3726 519216 3754
rect 513300 1222 513328 3726
rect 513288 1216 513340 1222
rect 513288 1158 513340 1164
rect 512184 1148 512236 1154
rect 512184 1090 512236 1096
rect 514496 1086 514524 3726
rect 514484 1080 514536 1086
rect 514484 1022 514536 1028
rect 510038 354 510150 480
rect 509712 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512430 82 512542 480
rect 513380 468 513432 474
rect 513380 410 513432 416
rect 513392 354 513420 410
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512104 66 512542 82
rect 512092 60 512542 66
rect 512144 54 512542 60
rect 512092 2 512144 8
rect 512430 -960 512542 54
rect 513534 -960 513646 326
rect 514730 218 514842 480
rect 514944 264 514996 270
rect 514730 212 514944 218
rect 514730 206 514996 212
rect 514730 190 514984 206
rect 514730 -960 514842 190
rect 515692 134 515720 3726
rect 515772 1352 515824 1358
rect 515772 1294 515824 1300
rect 515784 354 515812 1294
rect 515926 354 516038 480
rect 515784 326 516038 354
rect 515680 128 515732 134
rect 515680 70 515732 76
rect 515926 -960 516038 326
rect 516796 66 516824 3726
rect 517992 1290 518020 3726
rect 519188 1358 519216 3726
rect 520200 3726 520272 3754
rect 521440 3754 521468 4012
rect 522636 3754 522664 4012
rect 523740 3754 523768 4012
rect 524936 3754 524964 4012
rect 526040 3754 526068 4012
rect 527236 3754 527264 4012
rect 528432 3754 528460 4012
rect 529536 3754 529564 4012
rect 530732 3754 530760 4012
rect 531836 3754 531864 4012
rect 533032 3754 533060 4012
rect 534228 3754 534256 4012
rect 535332 3754 535360 4012
rect 536528 3754 536556 4012
rect 537632 3754 537660 4012
rect 538828 3754 538856 4012
rect 540024 3754 540052 4012
rect 541128 3754 541156 4012
rect 542324 3754 542352 4012
rect 521440 3726 521516 3754
rect 522636 3726 522712 3754
rect 523740 3726 523816 3754
rect 524936 3726 525012 3754
rect 526040 3726 526116 3754
rect 527236 3726 527312 3754
rect 528432 3726 528508 3754
rect 529536 3726 529612 3754
rect 530732 3726 530808 3754
rect 531836 3726 531912 3754
rect 533032 3726 533108 3754
rect 534228 3726 534304 3754
rect 535332 3726 535408 3754
rect 536528 3726 536604 3754
rect 537632 3726 537708 3754
rect 538828 3726 538904 3754
rect 540024 3726 540100 3754
rect 541128 3726 541204 3754
rect 519176 1352 519228 1358
rect 519176 1294 519228 1300
rect 517152 1284 517204 1290
rect 517152 1226 517204 1232
rect 517980 1284 518032 1290
rect 517980 1226 518032 1232
rect 517164 480 517192 1226
rect 519544 1216 519596 1222
rect 519544 1158 519596 1164
rect 517980 1148 518032 1154
rect 517980 1090 518032 1096
rect 516784 60 516836 66
rect 516784 2 516836 8
rect 517122 -960 517234 480
rect 517992 354 518020 1090
rect 519556 480 519584 1158
rect 520200 1018 520228 3726
rect 521488 1086 521516 3726
rect 522684 1222 522712 3726
rect 522672 1216 522724 1222
rect 522672 1158 522724 1164
rect 523788 1154 523816 3726
rect 523868 1284 523920 1290
rect 523868 1226 523920 1232
rect 523776 1148 523828 1154
rect 523776 1090 523828 1096
rect 520740 1080 520792 1086
rect 520740 1022 520792 1028
rect 521476 1080 521528 1086
rect 521476 1022 521528 1028
rect 520188 1012 520240 1018
rect 520188 954 520240 960
rect 520752 480 520780 1022
rect 518318 354 518430 480
rect 517992 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521660 128 521712 134
rect 521814 82 521926 480
rect 521712 76 521926 82
rect 521660 70 521926 76
rect 521672 54 521926 70
rect 521814 -960 521926 54
rect 523010 82 523122 480
rect 523880 354 523908 1226
rect 524206 354 524318 480
rect 523880 326 524318 354
rect 523010 66 523264 82
rect 523010 60 523276 66
rect 523010 54 523224 60
rect 523010 -960 523122 54
rect 523224 2 523276 8
rect 524206 -960 524318 326
rect 524984 134 525012 3726
rect 526088 1358 526116 3726
rect 525432 1352 525484 1358
rect 525432 1294 525484 1300
rect 526076 1352 526128 1358
rect 526076 1294 526128 1300
rect 525444 480 525472 1294
rect 527284 1290 527312 3726
rect 527272 1284 527324 1290
rect 527272 1226 527324 1232
rect 527824 1080 527876 1086
rect 527824 1022 527876 1028
rect 526628 1012 526680 1018
rect 526628 954 526680 960
rect 526640 480 526668 954
rect 527836 480 527864 1022
rect 524972 128 525024 134
rect 524972 70 525024 76
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528480 270 528508 3726
rect 529020 1216 529072 1222
rect 529020 1158 529072 1164
rect 529032 480 529060 1158
rect 529584 1086 529612 3726
rect 530780 1154 530808 3726
rect 531884 1222 531912 3726
rect 532148 1352 532200 1358
rect 532148 1294 532200 1300
rect 531872 1216 531924 1222
rect 531872 1158 531924 1164
rect 530124 1148 530176 1154
rect 530124 1090 530176 1096
rect 530768 1148 530820 1154
rect 530768 1090 530820 1096
rect 529572 1080 529624 1086
rect 529572 1022 529624 1028
rect 530136 480 530164 1090
rect 528468 264 528520 270
rect 528468 206 528520 212
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 82 531402 480
rect 532160 354 532188 1294
rect 533080 1018 533108 3726
rect 534276 1358 534304 3726
rect 534264 1352 534316 1358
rect 534264 1294 534316 1300
rect 533712 1284 533764 1290
rect 533712 1226 533764 1232
rect 533068 1012 533120 1018
rect 533068 954 533120 960
rect 533724 480 533752 1226
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 531504 128 531556 134
rect 531290 76 531504 82
rect 531290 70 531556 76
rect 531290 54 531544 70
rect 531290 -960 531402 54
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534540 264 534592 270
rect 534878 218 534990 480
rect 535380 406 535408 3726
rect 536104 1080 536156 1086
rect 536104 1022 536156 1028
rect 536116 480 536144 1022
rect 535368 400 535420 406
rect 535368 342 535420 348
rect 534592 212 534990 218
rect 534540 206 534990 212
rect 534552 190 534990 206
rect 534878 -960 534990 190
rect 536074 -960 536186 480
rect 536576 474 536604 3726
rect 537208 1148 537260 1154
rect 537208 1090 537260 1096
rect 537220 480 537248 1090
rect 536564 468 536616 474
rect 536564 410 536616 416
rect 537178 -960 537290 480
rect 537680 338 537708 3726
rect 538404 1216 538456 1222
rect 538404 1158 538456 1164
rect 538416 480 538444 1158
rect 538876 1154 538904 3726
rect 540072 1222 540100 3726
rect 540428 1352 540480 1358
rect 540428 1294 540480 1300
rect 540060 1216 540112 1222
rect 540060 1158 540112 1164
rect 538864 1148 538916 1154
rect 538864 1090 538916 1096
rect 539600 1012 539652 1018
rect 539600 954 539652 960
rect 539612 480 539640 954
rect 537668 332 537720 338
rect 537668 274 537720 280
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540440 354 540468 1294
rect 541176 746 541204 3726
rect 542280 3726 542352 3754
rect 543428 3754 543456 4012
rect 544624 3754 544652 4012
rect 545820 3754 545848 4012
rect 546924 3754 546952 4012
rect 548120 3754 548148 4012
rect 549316 3754 549344 4012
rect 550420 3754 550448 4012
rect 551616 3754 551644 4012
rect 552720 3754 552748 4012
rect 553916 3754 553944 4012
rect 555112 3754 555140 4012
rect 556216 3754 556244 4012
rect 557412 3754 557440 4012
rect 558516 3754 558544 4012
rect 559712 3754 559740 4012
rect 543428 3726 543504 3754
rect 544624 3726 544700 3754
rect 545820 3726 545896 3754
rect 546924 3726 547000 3754
rect 548120 3726 548196 3754
rect 549316 3726 549392 3754
rect 550420 3726 550496 3754
rect 551616 3726 551692 3754
rect 552720 3726 552796 3754
rect 553916 3726 553992 3754
rect 555112 3726 555188 3754
rect 556216 3726 556292 3754
rect 557412 3726 557488 3754
rect 542280 1358 542308 3726
rect 542268 1352 542320 1358
rect 542268 1294 542320 1300
rect 543476 1290 543504 3726
rect 543464 1284 543516 1290
rect 543464 1226 543516 1232
rect 541164 740 541216 746
rect 541164 682 541216 688
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 354 542074 480
rect 542820 468 542872 474
rect 542820 410 542872 416
rect 542176 400 542228 406
rect 541962 348 542176 354
rect 541962 342 542228 348
rect 542832 354 542860 410
rect 543158 354 543270 480
rect 541962 326 542216 342
rect 542832 326 543270 354
rect 541962 -960 542074 326
rect 543158 -960 543270 326
rect 544354 354 544466 480
rect 544672 474 544700 3726
rect 545488 1148 545540 1154
rect 545488 1090 545540 1096
rect 545500 480 545528 1090
rect 544660 468 544712 474
rect 544660 410 544712 416
rect 544354 338 544608 354
rect 544354 332 544620 338
rect 544354 326 544568 332
rect 544354 -960 544466 326
rect 544568 274 544620 280
rect 545458 -960 545570 480
rect 545868 338 545896 3726
rect 546684 1216 546736 1222
rect 546684 1158 546736 1164
rect 546696 480 546724 1158
rect 545856 332 545908 338
rect 545856 274 545908 280
rect 546654 -960 546766 480
rect 546972 406 547000 3726
rect 548168 1222 548196 3726
rect 549076 1352 549128 1358
rect 549076 1294 549128 1300
rect 548156 1216 548208 1222
rect 548156 1158 548208 1164
rect 547880 740 547932 746
rect 547880 682 547932 688
rect 547892 480 547920 682
rect 549088 480 549116 1294
rect 549364 1086 549392 3726
rect 550468 1290 550496 3726
rect 551664 1358 551692 3726
rect 551652 1352 551704 1358
rect 551652 1294 551704 1300
rect 550272 1284 550324 1290
rect 550272 1226 550324 1232
rect 550456 1284 550508 1290
rect 550456 1226 550508 1232
rect 549352 1080 549404 1086
rect 549352 1022 549404 1028
rect 550284 480 550312 1226
rect 552768 1154 552796 3726
rect 552756 1148 552808 1154
rect 552756 1090 552808 1096
rect 553964 678 553992 3726
rect 554964 1216 555016 1222
rect 554964 1158 555016 1164
rect 553952 672 554004 678
rect 552400 598 552704 626
rect 553952 614 554004 620
rect 546960 400 547012 406
rect 546960 342 547012 348
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551100 468 551152 474
rect 551100 410 551152 416
rect 551112 354 551140 410
rect 551438 354 551550 480
rect 551112 326 551550 354
rect 552400 338 552428 598
rect 552676 480 552704 598
rect 554976 480 555004 1158
rect 551438 -960 551550 326
rect 552388 332 552440 338
rect 552388 274 552440 280
rect 552634 -960 552746 480
rect 553738 354 553850 480
rect 553952 400 554004 406
rect 553738 348 553952 354
rect 553738 342 554004 348
rect 553738 326 553992 342
rect 553738 -960 553850 326
rect 554934 -960 555046 480
rect 555160 134 555188 3726
rect 556160 1080 556212 1086
rect 556160 1022 556212 1028
rect 556172 480 556200 1022
rect 556264 610 556292 3726
rect 557356 1284 557408 1290
rect 557356 1226 557408 1232
rect 556252 604 556304 610
rect 556252 546 556304 552
rect 557368 480 557396 1226
rect 557460 626 557488 3726
rect 558472 3726 558544 3754
rect 559668 3726 559740 3754
rect 560908 3754 560936 4012
rect 562012 3754 562040 4012
rect 563208 3754 563236 4012
rect 564312 3754 564340 4012
rect 565508 3754 565536 4012
rect 566704 3754 566732 4012
rect 560908 3726 560984 3754
rect 562012 3726 562088 3754
rect 558472 1222 558500 3726
rect 558552 1352 558604 1358
rect 558552 1294 558604 1300
rect 558460 1216 558512 1222
rect 558460 1158 558512 1164
rect 557540 740 557592 746
rect 557540 682 557592 688
rect 557552 626 557580 682
rect 557460 598 557580 626
rect 558564 480 558592 1294
rect 559668 1086 559696 3726
rect 560956 1358 560984 3726
rect 560944 1352 560996 1358
rect 560944 1294 560996 1300
rect 562060 1290 562088 3726
rect 563164 3726 563236 3754
rect 564268 3726 564340 3754
rect 565464 3726 565536 3754
rect 566660 3726 566732 3754
rect 567808 3754 567836 4012
rect 569004 3754 569032 4012
rect 570108 3754 570136 4012
rect 571304 3754 571332 4012
rect 567808 3726 567884 3754
rect 569004 3726 569080 3754
rect 570108 3726 570184 3754
rect 562048 1284 562100 1290
rect 562048 1226 562100 1232
rect 559748 1148 559800 1154
rect 559748 1090 559800 1096
rect 559656 1080 559708 1086
rect 559656 1022 559708 1028
rect 559760 480 559788 1090
rect 563164 678 563192 3726
rect 563152 672 563204 678
rect 563152 614 563204 620
rect 560852 604 560904 610
rect 560852 546 560904 552
rect 563244 604 563296 610
rect 563244 546 563296 552
rect 560864 480 560892 546
rect 563256 480 563284 546
rect 555148 128 555200 134
rect 555148 70 555200 76
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 82 562130 480
rect 562232 128 562284 134
rect 562018 76 562232 82
rect 562018 70 562284 76
rect 562018 54 562272 70
rect 562018 -960 562130 54
rect 563214 -960 563326 480
rect 564268 202 564296 3726
rect 564440 740 564492 746
rect 564440 682 564492 688
rect 564452 480 564480 682
rect 564256 196 564308 202
rect 564256 138 564308 144
rect 564410 -960 564522 480
rect 565464 134 565492 3726
rect 565636 1216 565688 1222
rect 565636 1158 565688 1164
rect 565648 480 565676 1158
rect 565452 128 565504 134
rect 565452 70 565504 76
rect 565606 -960 565718 480
rect 566660 474 566688 3726
rect 567856 1154 567884 3726
rect 568028 1352 568080 1358
rect 568028 1294 568080 1300
rect 567844 1148 567896 1154
rect 567844 1090 567896 1096
rect 566832 1080 566884 1086
rect 566832 1022 566884 1028
rect 566844 480 566872 1022
rect 568040 480 568068 1294
rect 569052 1222 569080 3726
rect 570156 1290 570184 3726
rect 571260 3726 571332 3754
rect 572500 3754 572528 4012
rect 573604 3754 573632 4012
rect 574800 3754 574828 4012
rect 575918 3998 576164 4026
rect 572500 3726 572576 3754
rect 573604 3726 573680 3754
rect 574800 3726 574876 3754
rect 571260 1358 571288 3726
rect 571248 1352 571300 1358
rect 571248 1294 571300 1300
rect 569132 1284 569184 1290
rect 569132 1226 569184 1232
rect 570144 1284 570196 1290
rect 570144 1226 570196 1232
rect 569040 1216 569092 1222
rect 569040 1158 569092 1164
rect 569144 480 569172 1226
rect 570328 672 570380 678
rect 570328 614 570380 620
rect 570340 480 570368 614
rect 566648 468 566700 474
rect 566648 410 566700 416
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 218 571606 480
rect 571352 202 571606 218
rect 571340 196 571606 202
rect 571392 190 571606 196
rect 571340 138 571392 144
rect 571494 -960 571606 190
rect 572548 66 572576 3726
rect 572690 82 572802 480
rect 573652 338 573680 3726
rect 573732 468 573784 474
rect 573732 410 573784 416
rect 573744 354 573772 410
rect 573886 354 573998 480
rect 573640 332 573692 338
rect 573744 326 573998 354
rect 573640 274 573692 280
rect 572904 128 572956 134
rect 572690 76 572904 82
rect 572690 70 572956 76
rect 572536 60 572588 66
rect 572536 2 572588 8
rect 572690 54 572944 70
rect 572690 -960 572802 54
rect 573886 -960 573998 326
rect 574848 202 574876 3726
rect 575112 1148 575164 1154
rect 575112 1090 575164 1096
rect 575124 480 575152 1090
rect 574836 196 574888 202
rect 574836 138 574888 144
rect 575082 -960 575194 480
rect 576136 134 576164 3998
rect 578608 1352 578660 1358
rect 578608 1294 578660 1300
rect 577412 1284 577464 1290
rect 577412 1226 577464 1232
rect 576308 1216 576360 1222
rect 576308 1158 576360 1164
rect 576320 480 576348 1158
rect 577424 480 577452 1226
rect 578620 480 578648 1294
rect 576124 128 576176 134
rect 576124 70 576176 76
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 82 579886 480
rect 579632 66 579886 82
rect 579620 60 579886 66
rect 579672 54 579886 60
rect 579620 2 579672 8
rect 579774 -960 579886 54
rect 580970 354 581082 480
rect 580970 338 581224 354
rect 580970 332 581236 338
rect 580970 326 581184 332
rect 580970 -960 581082 326
rect 581184 274 581236 280
rect 582166 218 582278 480
rect 581840 202 582278 218
rect 581828 196 582278 202
rect 581880 190 582278 196
rect 581828 138 581880 144
rect 582166 -960 582278 190
rect 583362 82 583474 480
rect 583576 128 583628 134
rect 583362 76 583576 82
rect 583362 70 583628 76
rect 583362 54 583616 70
rect 583362 -960 583474 54
<< via2 >>
rect 3514 697920 3570 697976
rect 576766 698128 576822 698184
rect 3514 697312 3570 697368
rect 580170 697176 580226 697232
rect 579526 684664 579582 684720
rect 579618 683848 579674 683904
rect 578330 644564 578386 644600
rect 578330 644544 578332 644564
rect 578332 644544 578384 644564
rect 578384 644544 578386 644564
rect 580906 644000 580962 644056
rect 3422 436600 3478 436656
rect 3422 435986 3478 436042
rect 3422 423544 3478 423600
rect 3422 422932 3478 422988
rect 3422 410488 3478 410544
rect 3422 409878 3478 409934
rect 3422 397432 3478 397488
rect 3422 396824 3478 396880
rect 3422 384376 3478 384432
rect 3422 383648 3478 383704
rect 3422 371320 3478 371376
rect 3422 370594 3478 370650
rect 3422 358400 3478 358456
rect 3422 357540 3478 357596
rect 579526 351872 579582 351928
rect 579526 351056 579582 351112
rect 3422 345344 3478 345400
rect 3422 344364 3478 344420
rect 579618 338544 579674 338600
rect 579526 337864 579582 337920
rect 3422 332288 3478 332344
rect 3422 331310 3478 331366
rect 580170 325216 580226 325272
rect 580170 324400 580226 324456
rect 3422 319232 3478 319288
rect 3422 318256 3478 318312
rect 579618 312024 579674 312080
rect 579526 311072 579582 311128
rect 3422 306176 3478 306232
rect 3422 305080 3478 305136
rect 579618 298696 579674 298752
rect 579526 297744 579582 297800
rect 3422 293120 3478 293176
rect 3422 292026 3478 292082
rect 580170 285368 580226 285424
rect 580170 284416 580226 284472
rect 3422 280064 3478 280120
rect 3422 278972 3478 279028
rect 579618 272176 579674 272232
rect 579526 271088 579582 271144
rect 3422 267144 3478 267200
rect 3422 265918 3478 265974
rect 580906 258848 580962 258904
rect 578882 257624 578938 257680
rect 3422 254088 3478 254144
rect 3422 252742 3478 252798
rect 580170 245520 580226 245576
rect 580170 244432 580226 244488
rect 3422 241032 3478 241088
rect 3422 239688 3478 239744
rect 579618 232328 579674 232384
rect 579526 231104 579582 231160
rect 3422 227976 3478 228032
rect 3422 226634 3478 226690
rect 579618 219000 579674 219056
rect 579526 217640 579582 217696
rect 3422 214920 3478 214976
rect 3422 213458 3478 213514
rect 579618 205672 579674 205728
rect 579526 204312 579582 204368
rect 3422 201864 3478 201920
rect 3422 200404 3478 200460
rect 579618 192480 579674 192536
rect 579526 190984 579582 191040
rect 3606 188808 3662 188864
rect 3606 187350 3662 187406
rect 579618 179152 579674 179208
rect 579526 177656 579582 177712
rect 3422 175888 3478 175944
rect 3422 174174 3478 174230
rect 579618 165824 579674 165880
rect 579526 164328 579582 164384
rect 2134 162832 2190 162888
rect 2134 161064 2190 161120
rect 580906 152632 580962 152688
rect 578514 151000 578570 151056
rect 3422 149776 3478 149832
rect 3422 148066 3478 148122
rect 579618 139304 579674 139360
rect 579526 137536 579582 137592
rect 2134 136720 2190 136776
rect 2134 134952 2190 135008
rect 579618 125976 579674 126032
rect 579526 124344 579582 124400
rect 3422 123664 3478 123720
rect 3422 121836 3478 121892
rect 579618 112784 579674 112840
rect 579526 110880 579582 110936
rect 2134 110608 2190 110664
rect 2134 108840 2190 108896
rect 579618 99456 579674 99512
rect 3422 97552 3478 97608
rect 579526 97552 579582 97608
rect 3422 95728 3478 95784
rect 579618 86128 579674 86184
rect 2134 84632 2190 84688
rect 579526 84224 579582 84280
rect 2134 82592 2190 82648
rect 579618 72936 579674 72992
rect 3422 71576 3478 71632
rect 579526 70896 579582 70952
rect 3422 69498 3478 69554
rect 579618 59608 579674 59664
rect 2134 58520 2190 58576
rect 579526 57568 579582 57624
rect 2134 56480 2190 56536
rect 579986 46280 580042 46336
rect 3422 45464 3478 45520
rect 578330 44240 578386 44296
rect 3422 43268 3478 43324
rect 579618 33088 579674 33144
rect 2134 32408 2190 32464
rect 579526 30912 579582 30968
rect 2134 30232 2190 30288
rect 579618 19760 579674 19816
rect 2042 19352 2098 19408
rect 579526 17584 579582 17640
rect 2042 17176 2098 17232
rect 579618 6568 579674 6624
rect 2778 6432 2834 6488
rect 2778 4120 2834 4176
rect 576766 4120 576822 4176
<< metal3 >>
rect 576761 698186 576827 698189
rect 575890 698184 576827 698186
rect 575890 698128 576766 698184
rect 576822 698128 576827 698184
rect 575890 698126 576827 698128
rect 3509 697978 3575 697981
rect 3509 697976 4048 697978
rect 3509 697920 3514 697976
rect 3570 697920 4048 697976
rect 575890 697948 575950 698126
rect 576761 698123 576827 698126
rect 3509 697918 4048 697920
rect 3509 697915 3575 697918
rect -960 697370 480 697460
rect 3509 697370 3575 697373
rect -960 697368 3575 697370
rect -960 697312 3514 697368
rect 3570 697312 3575 697368
rect -960 697310 3575 697312
rect -960 697220 480 697310
rect 3509 697307 3575 697310
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect 3374 684742 4048 684802
rect -960 684314 480 684404
rect 3374 684314 3434 684742
rect 579521 684722 579587 684725
rect 576350 684720 579587 684722
rect 576350 684680 579526 684720
rect 575920 684664 579526 684680
rect 579582 684664 579587 684720
rect 575920 684662 579587 684664
rect 575920 684620 576410 684662
rect 579521 684659 579587 684662
rect -960 684254 3434 684314
rect -960 684164 480 684254
rect 579613 683906 579679 683909
rect 583520 683906 584960 683996
rect 579613 683904 584960 683906
rect 579613 683848 579618 683904
rect 579674 683848 584960 683904
rect 579613 683846 584960 683848
rect 579613 683843 579679 683846
rect 583520 683756 584960 683846
rect 3374 671688 4048 671748
rect -960 671258 480 671348
rect 3374 671258 3434 671688
rect 576350 671382 583586 671394
rect 575920 671334 583586 671382
rect 575920 671322 576410 671334
rect -960 671198 3434 671258
rect -960 671108 480 671198
rect 583526 670850 583586 671334
rect 583342 670804 583586 670850
rect 583342 670790 584960 670804
rect 583342 670714 583402 670790
rect 583520 670714 584960 670790
rect 583342 670654 584960 670714
rect 583520 670564 584960 670654
rect 3374 658634 4048 658694
rect -960 658202 480 658292
rect 3374 658202 3434 658634
rect -960 658142 3434 658202
rect -960 658052 480 658142
rect 575920 657930 576410 657962
rect 575920 657902 583586 657930
rect 576350 657870 583586 657902
rect 583526 657522 583586 657870
rect 583342 657476 583586 657522
rect 583342 657462 584960 657476
rect 583342 657386 583402 657462
rect 583520 657386 584960 657462
rect 583342 657326 584960 657386
rect 583520 657236 584960 657326
rect 3374 645458 4048 645518
rect -960 645146 480 645236
rect 3374 645146 3434 645458
rect -960 645086 3434 645146
rect -960 644996 480 645086
rect 575920 644604 576410 644664
rect 576350 644602 576410 644604
rect 578325 644602 578391 644605
rect 576350 644600 578391 644602
rect 576350 644544 578330 644600
rect 578386 644544 578391 644600
rect 576350 644542 578391 644544
rect 578325 644539 578391 644542
rect 580901 644058 580967 644061
rect 583520 644058 584960 644148
rect 580901 644056 584960 644058
rect 580901 644000 580906 644056
rect 580962 644000 584960 644056
rect 580901 643998 584960 644000
rect 580901 643995 580967 643998
rect 583520 643908 584960 643998
rect 3374 632404 4048 632464
rect -960 632090 480 632180
rect 3374 632090 3434 632404
rect -960 632030 3434 632090
rect -960 631940 480 632030
rect 575920 631306 576410 631366
rect 576350 631274 576410 631306
rect 576350 631214 583586 631274
rect 583526 631002 583586 631214
rect 583342 630956 583586 631002
rect 583342 630942 584960 630956
rect 583342 630866 583402 630942
rect 583520 630866 584960 630942
rect 583342 630806 584960 630866
rect 583520 630716 584960 630806
rect 3374 619350 4048 619410
rect -960 619170 480 619260
rect 3374 619170 3434 619350
rect -960 619110 3434 619170
rect -960 619020 480 619110
rect 575920 617886 583586 617946
rect 583526 617674 583586 617886
rect 583342 617628 583586 617674
rect 583342 617614 584960 617628
rect 583342 617538 583402 617614
rect 583520 617538 584960 617614
rect 583342 617478 584960 617538
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3374 606174 4048 606234
rect 3374 606114 3434 606174
rect -960 606054 3434 606114
rect -960 605964 480 606054
rect 575920 604618 576410 604648
rect 575920 604588 576870 604618
rect 576350 604558 576870 604588
rect 576810 604482 576870 604558
rect 576810 604422 579722 604482
rect 579662 604210 579722 604422
rect 583520 604210 584960 604300
rect 579662 604150 584960 604210
rect 583520 604060 584960 604150
rect -960 593058 480 593148
rect 3374 593120 4048 593180
rect 3374 593058 3434 593120
rect -960 592998 3434 593058
rect -960 592908 480 592998
rect 575920 591290 576410 591350
rect 576350 591230 576870 591290
rect 576810 591018 576870 591230
rect 583520 591018 584960 591108
rect 576810 590958 584960 591018
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3374 580066 4048 580126
rect 3374 580002 3434 580066
rect -960 579942 3434 580002
rect -960 579852 480 579942
rect 575920 577870 576410 577930
rect 576350 577826 576410 577870
rect 576350 577766 576870 577826
rect 576810 577690 576870 577766
rect 583520 577690 584960 577780
rect 576810 577630 584960 577690
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3374 566946 4048 566950
rect -960 566890 4048 566946
rect -960 566886 3434 566890
rect -960 566796 480 566886
rect 575920 564572 576410 564632
rect 576350 564498 576410 564572
rect 576350 564438 579722 564498
rect 579662 564362 579722 564438
rect 583520 564362 584960 564452
rect 579662 564302 584960 564362
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3374 553890 4048 553896
rect -960 553836 4048 553890
rect -960 553830 3434 553836
rect -960 553740 480 553830
rect 575920 551170 576410 551212
rect 583520 551170 584960 551260
rect 575920 551152 584960 551170
rect 576350 551110 584960 551152
rect 583520 551020 584960 551110
rect -960 540834 480 540924
rect 3374 540834 4048 540842
rect -960 540782 4048 540834
rect -960 540774 3434 540782
rect -960 540684 480 540774
rect 575920 537854 576410 537914
rect 576350 537842 576410 537854
rect 583520 537842 584960 537932
rect 576350 537782 584960 537842
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect -960 527854 3434 527914
rect -960 527764 480 527854
rect 3374 527788 3434 527854
rect 3374 527728 4048 527788
rect 575920 524556 576410 524616
rect 576350 524514 576410 524556
rect 583520 524514 584960 524604
rect 576350 524454 584960 524514
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect -960 514798 3434 514858
rect -960 514708 480 514798
rect 3374 514612 3434 514798
rect 3374 514552 4048 514612
rect 583520 511322 584960 511412
rect 576350 511262 584960 511322
rect 576350 511196 576410 511262
rect 575920 511136 576410 511196
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect -960 501742 3434 501802
rect -960 501652 480 501742
rect 3374 501558 3434 501742
rect 3374 501498 4048 501558
rect 583520 497994 584960 498084
rect 576350 497934 584960 497994
rect 576350 497898 576410 497934
rect 575920 497838 576410 497898
rect 583520 497844 584960 497934
rect -960 488746 480 488836
rect -960 488686 3434 488746
rect -960 488596 480 488686
rect 3374 488504 3434 488686
rect 3374 488444 4048 488504
rect 583520 484666 584960 484756
rect 576350 484606 584960 484666
rect 576350 484600 576410 484606
rect 575920 484540 576410 484600
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect -960 475630 3434 475690
rect -960 475540 480 475630
rect 3374 475328 3434 475630
rect 3374 475268 4048 475328
rect 583520 471474 584960 471564
rect 576810 471414 584960 471474
rect 576810 471202 576870 471414
rect 583520 471324 584960 471414
rect 576350 471180 576870 471202
rect 575920 471142 576870 471180
rect 575920 471120 576410 471142
rect -960 462634 480 462724
rect -960 462574 3434 462634
rect -960 462484 480 462574
rect 3374 462274 3434 462574
rect 3374 462214 4048 462274
rect 583520 458146 584960 458236
rect 576810 458086 584960 458146
rect 576810 458010 576870 458086
rect 576350 457950 576870 458010
rect 583520 457996 584960 458086
rect 576350 457882 576410 457950
rect 575920 457822 576410 457882
rect -960 449578 480 449668
rect -960 449518 3434 449578
rect -960 449428 480 449518
rect 3374 449220 3434 449518
rect 3374 449160 4048 449220
rect 583520 444818 584960 444908
rect 576810 444758 584960 444818
rect 576810 444682 576870 444758
rect 576350 444622 576870 444682
rect 583520 444668 584960 444758
rect 576350 444584 576410 444622
rect 575920 444524 576410 444584
rect -960 436658 480 436748
rect 3417 436658 3483 436661
rect -960 436656 3483 436658
rect -960 436600 3422 436656
rect 3478 436600 3483 436656
rect -960 436598 3483 436600
rect -960 436508 480 436598
rect 3417 436595 3483 436598
rect 3417 436044 3483 436047
rect 3417 436042 4048 436044
rect 3417 435986 3422 436042
rect 3478 435986 4048 436042
rect 3417 435984 4048 435986
rect 3417 435981 3483 435984
rect 583520 431626 584960 431716
rect 583342 431566 584960 431626
rect 583342 431490 583402 431566
rect 583520 431490 584960 431566
rect 583342 431476 584960 431490
rect 583342 431430 583586 431476
rect 583526 431218 583586 431430
rect 576350 431164 583586 431218
rect 575920 431158 583586 431164
rect 575920 431104 576410 431158
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 3417 422990 3483 422993
rect 3417 422988 4048 422990
rect 3417 422932 3422 422988
rect 3478 422932 4048 422988
rect 3417 422930 4048 422932
rect 3417 422927 3483 422930
rect 583520 418298 584960 418388
rect 579662 418238 584960 418298
rect 579662 418162 579722 418238
rect 576810 418102 579722 418162
rect 583520 418148 584960 418238
rect 576810 417890 576870 418102
rect 576350 417866 576870 417890
rect 575920 417830 576870 417866
rect 575920 417806 576410 417830
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 3417 409936 3483 409939
rect 3417 409934 4048 409936
rect 3417 409878 3422 409934
rect 3478 409878 4048 409934
rect 3417 409876 4048 409878
rect 3417 409873 3483 409876
rect 583520 404970 584960 405060
rect 583342 404910 584960 404970
rect 583342 404834 583402 404910
rect 583520 404834 584960 404910
rect 583342 404820 584960 404834
rect 583342 404774 583586 404820
rect 583526 404562 583586 404774
rect 576350 404502 583586 404562
rect 576350 404446 576410 404502
rect 575920 404386 576410 404446
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 3417 396882 3483 396885
rect 3417 396880 4048 396882
rect 3417 396824 3422 396880
rect 3478 396824 4048 396880
rect 3417 396822 4048 396824
rect 3417 396819 3483 396822
rect 583520 391778 584960 391868
rect 583342 391718 584960 391778
rect 583342 391642 583402 391718
rect 583520 391642 584960 391718
rect 583342 391628 584960 391642
rect 583342 391582 583586 391628
rect 583526 391234 583586 391582
rect 576350 391174 583586 391234
rect 576350 391148 576410 391174
rect 575920 391088 576410 391148
rect -960 384434 480 384524
rect 3417 384434 3483 384437
rect -960 384432 3483 384434
rect -960 384376 3422 384432
rect 3478 384376 3483 384432
rect -960 384374 3483 384376
rect -960 384284 480 384374
rect 3417 384371 3483 384374
rect 3417 383706 3483 383709
rect 3417 383704 4048 383706
rect 3417 383648 3422 383704
rect 3478 383648 4048 383704
rect 3417 383646 4048 383648
rect 3417 383643 3483 383646
rect 583520 378450 584960 378540
rect 579662 378390 584960 378450
rect 579662 378178 579722 378390
rect 583520 378300 584960 378390
rect 579478 378118 579722 378178
rect 579478 377906 579538 378118
rect 576350 377850 579538 377906
rect 575920 377846 579538 377850
rect 575920 377790 576410 377846
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 3417 370652 3483 370655
rect 3417 370650 4048 370652
rect 3417 370594 3422 370650
rect 3478 370594 4048 370650
rect 3417 370592 4048 370594
rect 3417 370589 3483 370592
rect 583520 365122 584960 365212
rect 583342 365062 584960 365122
rect 583342 364986 583402 365062
rect 583520 364986 584960 365062
rect 583342 364972 584960 364986
rect 583342 364926 583586 364972
rect 583526 364442 583586 364926
rect 576350 364430 583586 364442
rect 575920 364382 583586 364430
rect 575920 364370 576410 364382
rect -960 358458 480 358548
rect 3417 358458 3483 358461
rect -960 358456 3483 358458
rect -960 358400 3422 358456
rect 3478 358400 3483 358456
rect -960 358398 3483 358400
rect -960 358308 480 358398
rect 3417 358395 3483 358398
rect 3417 357598 3483 357601
rect 3417 357596 4048 357598
rect 3417 357540 3422 357596
rect 3478 357540 4048 357596
rect 3417 357538 4048 357540
rect 3417 357535 3483 357538
rect 579521 351930 579587 351933
rect 583520 351930 584960 352020
rect 579521 351928 584960 351930
rect 579521 351872 579526 351928
rect 579582 351872 584960 351928
rect 579521 351870 584960 351872
rect 579521 351867 579587 351870
rect 583520 351780 584960 351870
rect 575920 351114 576410 351132
rect 579521 351114 579587 351117
rect 575920 351112 579587 351114
rect 575920 351072 579526 351112
rect 576350 351056 579526 351072
rect 579582 351056 579587 351112
rect 576350 351054 579587 351056
rect 579521 351051 579587 351054
rect -960 345402 480 345492
rect 3417 345402 3483 345405
rect -960 345400 3483 345402
rect -960 345344 3422 345400
rect 3478 345344 3483 345400
rect -960 345342 3483 345344
rect -960 345252 480 345342
rect 3417 345339 3483 345342
rect 3417 344422 3483 344425
rect 3417 344420 4048 344422
rect 3417 344364 3422 344420
rect 3478 344364 4048 344420
rect 3417 344362 4048 344364
rect 3417 344359 3483 344362
rect 579613 338602 579679 338605
rect 583520 338602 584960 338692
rect 579613 338600 584960 338602
rect 579613 338544 579618 338600
rect 579674 338544 584960 338600
rect 579613 338542 584960 338544
rect 579613 338539 579679 338542
rect 583520 338452 584960 338542
rect 579521 337922 579587 337925
rect 576350 337920 579587 337922
rect 576350 337864 579526 337920
rect 579582 337864 579587 337920
rect 576350 337862 579587 337864
rect 576350 337834 576410 337862
rect 579521 337859 579587 337862
rect 575920 337774 576410 337834
rect -960 332346 480 332436
rect 3417 332346 3483 332349
rect -960 332344 3483 332346
rect -960 332288 3422 332344
rect 3478 332288 3483 332344
rect -960 332286 3483 332288
rect -960 332196 480 332286
rect 3417 332283 3483 332286
rect 3417 331368 3483 331371
rect 3417 331366 4048 331368
rect 3417 331310 3422 331366
rect 3478 331310 4048 331366
rect 3417 331308 4048 331310
rect 3417 331305 3483 331308
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 580165 324458 580231 324461
rect 576350 324456 580231 324458
rect 576350 324414 580170 324456
rect 575920 324400 580170 324414
rect 580226 324400 580231 324456
rect 575920 324398 580231 324400
rect 575920 324354 576410 324398
rect 580165 324395 580231 324398
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 3417 318314 3483 318317
rect 3417 318312 4048 318314
rect 3417 318256 3422 318312
rect 3478 318256 4048 318312
rect 3417 318254 4048 318256
rect 3417 318251 3483 318254
rect 579613 312082 579679 312085
rect 583520 312082 584960 312172
rect 579613 312080 584960 312082
rect 579613 312024 579618 312080
rect 579674 312024 584960 312080
rect 579613 312022 584960 312024
rect 579613 312019 579679 312022
rect 583520 311932 584960 312022
rect 579521 311130 579587 311133
rect 576350 311128 579587 311130
rect 576350 311116 579526 311128
rect 575920 311072 579526 311116
rect 579582 311072 579587 311128
rect 575920 311070 579587 311072
rect 575920 311056 576410 311070
rect 579521 311067 579587 311070
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 3417 305138 3483 305141
rect 3417 305136 4048 305138
rect 3417 305080 3422 305136
rect 3478 305080 4048 305136
rect 3417 305078 4048 305080
rect 3417 305075 3483 305078
rect 579613 298754 579679 298757
rect 583520 298754 584960 298844
rect 579613 298752 584960 298754
rect 579613 298696 579618 298752
rect 579674 298696 584960 298752
rect 579613 298694 584960 298696
rect 579613 298691 579679 298694
rect 583520 298604 584960 298694
rect 575920 297802 576410 297818
rect 579521 297802 579587 297805
rect 575920 297800 579587 297802
rect 575920 297758 579526 297800
rect 576350 297744 579526 297758
rect 579582 297744 579587 297800
rect 576350 297742 579587 297744
rect 579521 297739 579587 297742
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 3417 292084 3483 292087
rect 3417 292082 4048 292084
rect 3417 292026 3422 292082
rect 3478 292026 4048 292082
rect 3417 292024 4048 292026
rect 3417 292021 3483 292024
rect 580165 285426 580231 285429
rect 583520 285426 584960 285516
rect 580165 285424 584960 285426
rect 580165 285368 580170 285424
rect 580226 285368 584960 285424
rect 580165 285366 584960 285368
rect 580165 285363 580231 285366
rect 583520 285276 584960 285366
rect 580165 284474 580231 284477
rect 576350 284472 580231 284474
rect 576350 284416 580170 284472
rect 580226 284416 580231 284472
rect 576350 284414 580231 284416
rect 576350 284398 576410 284414
rect 580165 284411 580231 284414
rect 575920 284338 576410 284398
rect -960 280122 480 280212
rect 3417 280122 3483 280125
rect -960 280120 3483 280122
rect -960 280064 3422 280120
rect 3478 280064 3483 280120
rect -960 280062 3483 280064
rect -960 279972 480 280062
rect 3417 280059 3483 280062
rect 3417 279030 3483 279033
rect 3417 279028 4048 279030
rect 3417 278972 3422 279028
rect 3478 278972 4048 279028
rect 3417 278970 4048 278972
rect 3417 278967 3483 278970
rect 579613 272234 579679 272237
rect 583520 272234 584960 272324
rect 579613 272232 584960 272234
rect 579613 272176 579618 272232
rect 579674 272176 584960 272232
rect 579613 272174 584960 272176
rect 579613 272171 579679 272174
rect 583520 272084 584960 272174
rect 579521 271146 579587 271149
rect 576350 271144 579587 271146
rect 576350 271100 579526 271144
rect 575920 271088 579526 271100
rect 579582 271088 579587 271144
rect 575920 271086 579587 271088
rect 575920 271040 576410 271086
rect 579521 271083 579587 271086
rect -960 267202 480 267292
rect 3417 267202 3483 267205
rect -960 267200 3483 267202
rect -960 267144 3422 267200
rect 3478 267144 3483 267200
rect -960 267142 3483 267144
rect -960 267052 480 267142
rect 3417 267139 3483 267142
rect 3417 265976 3483 265979
rect 3417 265974 4048 265976
rect 3417 265918 3422 265974
rect 3478 265918 4048 265974
rect 3417 265916 4048 265918
rect 3417 265913 3483 265916
rect 580901 258906 580967 258909
rect 583520 258906 584960 258996
rect 580901 258904 584960 258906
rect 580901 258848 580906 258904
rect 580962 258848 584960 258904
rect 580901 258846 584960 258848
rect 580901 258843 580967 258846
rect 583520 258756 584960 258846
rect 578877 257682 578943 257685
rect 576350 257680 578943 257682
rect 575920 257624 578882 257680
rect 578938 257624 578943 257680
rect 575920 257622 578943 257624
rect 575920 257620 576410 257622
rect 578877 257619 578943 257622
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 3417 252800 3483 252803
rect 3417 252798 4048 252800
rect 3417 252742 3422 252798
rect 3478 252742 4048 252798
rect 3417 252740 4048 252742
rect 3417 252737 3483 252740
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 580165 244490 580231 244493
rect 576350 244488 580231 244490
rect 576350 244432 580170 244488
rect 580226 244432 580231 244488
rect 576350 244430 580231 244432
rect 576350 244382 576410 244430
rect 580165 244427 580231 244430
rect 575920 244322 576410 244382
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 3417 239746 3483 239749
rect 3417 239744 4048 239746
rect 3417 239688 3422 239744
rect 3478 239688 4048 239744
rect 3417 239686 4048 239688
rect 3417 239683 3483 239686
rect 579613 232386 579679 232389
rect 583520 232386 584960 232476
rect 579613 232384 584960 232386
rect 579613 232328 579618 232384
rect 579674 232328 584960 232384
rect 579613 232326 584960 232328
rect 579613 232323 579679 232326
rect 583520 232236 584960 232326
rect 579521 231162 579587 231165
rect 576350 231160 579587 231162
rect 576350 231104 579526 231160
rect 579582 231104 579587 231160
rect 576350 231102 579587 231104
rect 576350 231084 576410 231102
rect 579521 231099 579587 231102
rect 575920 231024 576410 231084
rect -960 228034 480 228124
rect 3417 228034 3483 228037
rect -960 228032 3483 228034
rect -960 227976 3422 228032
rect 3478 227976 3483 228032
rect -960 227974 3483 227976
rect -960 227884 480 227974
rect 3417 227971 3483 227974
rect 3417 226692 3483 226695
rect 3417 226690 4048 226692
rect 3417 226634 3422 226690
rect 3478 226634 4048 226690
rect 3417 226632 4048 226634
rect 3417 226629 3483 226632
rect 579613 219058 579679 219061
rect 583520 219058 584960 219148
rect 579613 219056 584960 219058
rect 579613 219000 579618 219056
rect 579674 219000 584960 219056
rect 579613 218998 584960 219000
rect 579613 218995 579679 218998
rect 583520 218908 584960 218998
rect 579521 217698 579587 217701
rect 576350 217696 579587 217698
rect 576350 217664 579526 217696
rect 575920 217640 579526 217664
rect 579582 217640 579587 217696
rect 575920 217638 579587 217640
rect 575920 217604 576410 217638
rect 579521 217635 579587 217638
rect -960 214978 480 215068
rect 3417 214978 3483 214981
rect -960 214976 3483 214978
rect -960 214920 3422 214976
rect 3478 214920 3483 214976
rect -960 214918 3483 214920
rect -960 214828 480 214918
rect 3417 214915 3483 214918
rect 3417 213516 3483 213519
rect 3417 213514 4048 213516
rect 3417 213458 3422 213514
rect 3478 213458 4048 213514
rect 3417 213456 4048 213458
rect 3417 213453 3483 213456
rect 579613 205730 579679 205733
rect 583520 205730 584960 205820
rect 579613 205728 584960 205730
rect 579613 205672 579618 205728
rect 579674 205672 584960 205728
rect 579613 205670 584960 205672
rect 579613 205667 579679 205670
rect 583520 205580 584960 205670
rect 579521 204370 579587 204373
rect 576350 204368 579587 204370
rect 576350 204366 579526 204368
rect 575920 204312 579526 204366
rect 579582 204312 579587 204368
rect 575920 204310 579587 204312
rect 575920 204306 576410 204310
rect 579521 204307 579587 204310
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 3417 200462 3483 200465
rect 3417 200460 4048 200462
rect 3417 200404 3422 200460
rect 3478 200404 4048 200460
rect 3417 200402 4048 200404
rect 3417 200399 3483 200402
rect 579613 192538 579679 192541
rect 583520 192538 584960 192628
rect 579613 192536 584960 192538
rect 579613 192480 579618 192536
rect 579674 192480 584960 192536
rect 579613 192478 584960 192480
rect 579613 192475 579679 192478
rect 583520 192388 584960 192478
rect 575920 191042 576410 191068
rect 579521 191042 579587 191045
rect 575920 191040 579587 191042
rect 575920 191008 579526 191040
rect 576350 190984 579526 191008
rect 579582 190984 579587 191040
rect 576350 190982 579587 190984
rect 579521 190979 579587 190982
rect -960 188866 480 188956
rect 3601 188866 3667 188869
rect -960 188864 3667 188866
rect -960 188808 3606 188864
rect 3662 188808 3667 188864
rect -960 188806 3667 188808
rect -960 188716 480 188806
rect 3601 188803 3667 188806
rect 3601 187408 3667 187411
rect 3601 187406 4048 187408
rect 3601 187350 3606 187406
rect 3662 187350 4048 187406
rect 3601 187348 4048 187350
rect 3601 187345 3667 187348
rect 579613 179210 579679 179213
rect 583520 179210 584960 179300
rect 579613 179208 584960 179210
rect 579613 179152 579618 179208
rect 579674 179152 584960 179208
rect 579613 179150 584960 179152
rect 579613 179147 579679 179150
rect 583520 179060 584960 179150
rect 579521 177714 579587 177717
rect 576350 177712 579587 177714
rect 576350 177656 579526 177712
rect 579582 177656 579587 177712
rect 576350 177654 579587 177656
rect 576350 177648 576410 177654
rect 579521 177651 579587 177654
rect 575920 177588 576410 177648
rect -960 175946 480 176036
rect 3417 175946 3483 175949
rect -960 175944 3483 175946
rect -960 175888 3422 175944
rect 3478 175888 3483 175944
rect -960 175886 3483 175888
rect -960 175796 480 175886
rect 3417 175883 3483 175886
rect 3417 174232 3483 174235
rect 3417 174230 4048 174232
rect 3417 174174 3422 174230
rect 3478 174174 4048 174230
rect 3417 174172 4048 174174
rect 3417 174169 3483 174172
rect 579613 165882 579679 165885
rect 583520 165882 584960 165972
rect 579613 165880 584960 165882
rect 579613 165824 579618 165880
rect 579674 165824 584960 165880
rect 579613 165822 584960 165824
rect 579613 165819 579679 165822
rect 583520 165732 584960 165822
rect 579521 164386 579587 164389
rect 576350 164384 579587 164386
rect 576350 164350 579526 164384
rect 575920 164328 579526 164350
rect 579582 164328 579587 164384
rect 575920 164326 579587 164328
rect 575920 164290 576410 164326
rect 579521 164323 579587 164326
rect -960 162890 480 162980
rect 2129 162890 2195 162893
rect -960 162888 2195 162890
rect -960 162832 2134 162888
rect 2190 162832 2195 162888
rect -960 162830 2195 162832
rect -960 162740 480 162830
rect 2129 162827 2195 162830
rect 2129 161122 2195 161125
rect 3374 161122 4048 161178
rect 2129 161120 4048 161122
rect 2129 161064 2134 161120
rect 2190 161118 4048 161120
rect 2190 161064 3434 161118
rect 2129 161062 3434 161064
rect 2129 161059 2195 161062
rect 580901 152690 580967 152693
rect 583520 152690 584960 152780
rect 580901 152688 584960 152690
rect 580901 152632 580906 152688
rect 580962 152632 584960 152688
rect 580901 152630 584960 152632
rect 580901 152627 580967 152630
rect 583520 152540 584960 152630
rect 578509 151058 578575 151061
rect 576350 151056 578575 151058
rect 576350 151052 578514 151056
rect 575920 151000 578514 151052
rect 578570 151000 578575 151056
rect 575920 150998 578575 151000
rect 575920 150992 576410 150998
rect 578509 150995 578575 150998
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 3417 148124 3483 148127
rect 3417 148122 4048 148124
rect 3417 148066 3422 148122
rect 3478 148066 4048 148122
rect 3417 148064 4048 148066
rect 3417 148061 3483 148064
rect 579613 139362 579679 139365
rect 583520 139362 584960 139452
rect 579613 139360 584960 139362
rect 579613 139304 579618 139360
rect 579674 139304 584960 139360
rect 579613 139302 584960 139304
rect 579613 139299 579679 139302
rect 583520 139212 584960 139302
rect 575920 137594 576410 137632
rect 579521 137594 579587 137597
rect 575920 137592 579587 137594
rect 575920 137572 579526 137592
rect 576350 137536 579526 137572
rect 579582 137536 579587 137592
rect 576350 137534 579587 137536
rect 579521 137531 579587 137534
rect -960 136778 480 136868
rect 2129 136778 2195 136781
rect -960 136776 2195 136778
rect -960 136720 2134 136776
rect 2190 136720 2195 136776
rect -960 136718 2195 136720
rect -960 136628 480 136718
rect 2129 136715 2195 136718
rect 2129 135010 2195 135013
rect 3374 135010 4048 135070
rect 2129 135008 3434 135010
rect 2129 134952 2134 135008
rect 2190 134952 3434 135008
rect 2129 134950 3434 134952
rect 2129 134947 2195 134950
rect 579613 126034 579679 126037
rect 583520 126034 584960 126124
rect 579613 126032 584960 126034
rect 579613 125976 579618 126032
rect 579674 125976 584960 126032
rect 579613 125974 584960 125976
rect 579613 125971 579679 125974
rect 583520 125884 584960 125974
rect 579521 124402 579587 124405
rect 576350 124400 579587 124402
rect 576350 124344 579526 124400
rect 579582 124344 579587 124400
rect 576350 124342 579587 124344
rect 576350 124334 576410 124342
rect 579521 124339 579587 124342
rect 575920 124274 576410 124334
rect -960 123722 480 123812
rect 3417 123722 3483 123725
rect -960 123720 3483 123722
rect -960 123664 3422 123720
rect 3478 123664 3483 123720
rect -960 123662 3483 123664
rect -960 123572 480 123662
rect 3417 123659 3483 123662
rect 3417 121894 3483 121897
rect 3417 121892 4048 121894
rect 3417 121836 3422 121892
rect 3478 121836 4048 121892
rect 3417 121834 4048 121836
rect 3417 121831 3483 121834
rect 579613 112842 579679 112845
rect 583520 112842 584960 112932
rect 579613 112840 584960 112842
rect 579613 112784 579618 112840
rect 579674 112784 584960 112840
rect 579613 112782 584960 112784
rect 579613 112779 579679 112782
rect 583520 112692 584960 112782
rect 579521 110938 579587 110941
rect 576350 110936 579587 110938
rect 576350 110914 579526 110936
rect 575920 110880 579526 110914
rect 579582 110880 579587 110936
rect 575920 110878 579587 110880
rect 575920 110854 576410 110878
rect 579521 110875 579587 110878
rect -960 110666 480 110756
rect 2129 110666 2195 110669
rect -960 110664 2195 110666
rect -960 110608 2134 110664
rect 2190 110608 2195 110664
rect -960 110606 2195 110608
rect -960 110516 480 110606
rect 2129 110603 2195 110606
rect 2129 108898 2195 108901
rect 2129 108896 3434 108898
rect 2129 108840 2134 108896
rect 2190 108840 3434 108896
rect 2129 108838 4048 108840
rect 2129 108835 2195 108838
rect 3374 108780 4048 108838
rect 579613 99514 579679 99517
rect 583520 99514 584960 99604
rect 579613 99512 584960 99514
rect 579613 99456 579618 99512
rect 579674 99456 584960 99512
rect 579613 99454 584960 99456
rect 579613 99451 579679 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect 575920 97610 576410 97616
rect 579521 97610 579587 97613
rect 575920 97608 579587 97610
rect 575920 97556 579526 97608
rect -960 97550 3483 97552
rect 576350 97552 579526 97556
rect 579582 97552 579587 97608
rect 576350 97550 579587 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 579521 97547 579587 97550
rect 3417 95786 3483 95789
rect 3417 95784 4048 95786
rect 3417 95728 3422 95784
rect 3478 95728 4048 95784
rect 3417 95726 4048 95728
rect 3417 95723 3483 95726
rect 579613 86186 579679 86189
rect 583520 86186 584960 86276
rect 579613 86184 584960 86186
rect 579613 86128 579618 86184
rect 579674 86128 584960 86184
rect 579613 86126 584960 86128
rect 579613 86123 579679 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 2129 84690 2195 84693
rect -960 84688 2195 84690
rect -960 84632 2134 84688
rect 2190 84632 2195 84688
rect -960 84630 2195 84632
rect -960 84540 480 84630
rect 2129 84627 2195 84630
rect 575920 84282 576410 84318
rect 579521 84282 579587 84285
rect 575920 84280 579587 84282
rect 575920 84258 579526 84280
rect 576350 84224 579526 84258
rect 579582 84224 579587 84280
rect 576350 84222 579587 84224
rect 579521 84219 579587 84222
rect 2129 82650 2195 82653
rect 2129 82648 3434 82650
rect 2129 82592 2134 82648
rect 2190 82610 3434 82648
rect 2190 82592 4048 82610
rect 2129 82590 4048 82592
rect 2129 82587 2195 82590
rect 3374 82550 4048 82590
rect 579613 72994 579679 72997
rect 583520 72994 584960 73084
rect 579613 72992 584960 72994
rect 579613 72936 579618 72992
rect 579674 72936 584960 72992
rect 579613 72934 584960 72936
rect 579613 72931 579679 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 579521 70954 579587 70957
rect 576350 70952 579587 70954
rect 576350 70898 579526 70952
rect 575920 70896 579526 70898
rect 579582 70896 579587 70952
rect 575920 70894 579587 70896
rect 575920 70838 576410 70894
rect 579521 70891 579587 70894
rect 3417 69556 3483 69559
rect 3417 69554 4048 69556
rect 3417 69498 3422 69554
rect 3478 69498 4048 69554
rect 3417 69496 4048 69498
rect 3417 69493 3483 69496
rect 579613 59666 579679 59669
rect 583520 59666 584960 59756
rect 579613 59664 584960 59666
rect 579613 59608 579618 59664
rect 579674 59608 584960 59664
rect 579613 59606 584960 59608
rect 579613 59603 579679 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 2129 58578 2195 58581
rect -960 58576 2195 58578
rect -960 58520 2134 58576
rect 2190 58520 2195 58576
rect -960 58518 2195 58520
rect -960 58428 480 58518
rect 2129 58515 2195 58518
rect 579521 57626 579587 57629
rect 576350 57624 579587 57626
rect 576350 57600 579526 57624
rect 575920 57568 579526 57600
rect 579582 57568 579587 57624
rect 575920 57566 579587 57568
rect 575920 57540 576410 57566
rect 579521 57563 579587 57566
rect 2129 56538 2195 56541
rect 2129 56536 3434 56538
rect 2129 56480 2134 56536
rect 2190 56502 3434 56536
rect 2190 56480 4048 56502
rect 2129 56478 4048 56480
rect 2129 56475 2195 56478
rect 3374 56442 4048 56478
rect 579981 46338 580047 46341
rect 583520 46338 584960 46428
rect 579981 46336 584960 46338
rect 579981 46280 579986 46336
rect 580042 46280 584960 46336
rect 579981 46278 584960 46280
rect 579981 46275 580047 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 575920 44298 576410 44302
rect 578325 44298 578391 44301
rect 575920 44296 578391 44298
rect 575920 44242 578330 44296
rect 576350 44240 578330 44242
rect 578386 44240 578391 44296
rect 576350 44238 578391 44240
rect 578325 44235 578391 44238
rect 3417 43326 3483 43329
rect 3417 43324 4048 43326
rect 3417 43268 3422 43324
rect 3478 43268 4048 43324
rect 3417 43266 4048 43268
rect 3417 43263 3483 43266
rect 579613 33146 579679 33149
rect 583520 33146 584960 33236
rect 579613 33144 584960 33146
rect 579613 33088 579618 33144
rect 579674 33088 584960 33144
rect 579613 33086 584960 33088
rect 579613 33083 579679 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2129 32466 2195 32469
rect -960 32464 2195 32466
rect -960 32408 2134 32464
rect 2190 32408 2195 32464
rect -960 32406 2195 32408
rect -960 32316 480 32406
rect 2129 32403 2195 32406
rect 579521 30970 579587 30973
rect 576350 30968 579587 30970
rect 576350 30912 579526 30968
rect 579582 30912 579587 30968
rect 576350 30910 579587 30912
rect 576350 30882 576410 30910
rect 579521 30907 579587 30910
rect 575920 30822 576410 30882
rect 2129 30290 2195 30293
rect 2129 30288 3434 30290
rect 2129 30232 2134 30288
rect 2190 30272 3434 30288
rect 2190 30232 4048 30272
rect 2129 30230 4048 30232
rect 2129 30227 2195 30230
rect 3374 30212 4048 30230
rect 579613 19818 579679 19821
rect 583520 19818 584960 19908
rect 579613 19816 584960 19818
rect 579613 19760 579618 19816
rect 579674 19760 584960 19816
rect 579613 19758 584960 19760
rect 579613 19755 579679 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 2037 19410 2103 19413
rect -960 19408 2103 19410
rect -960 19352 2042 19408
rect 2098 19352 2103 19408
rect -960 19350 2103 19352
rect -960 19260 480 19350
rect 2037 19347 2103 19350
rect 579521 17642 579587 17645
rect 576350 17640 579587 17642
rect 576350 17584 579526 17640
rect 579582 17584 579587 17640
rect 575920 17582 579587 17584
rect 575920 17524 576410 17582
rect 579521 17579 579587 17582
rect 2037 17234 2103 17237
rect 2037 17232 3434 17234
rect 2037 17176 2042 17232
rect 2098 17218 3434 17232
rect 2098 17176 4048 17218
rect 2037 17174 4048 17176
rect 2037 17171 2103 17174
rect 3374 17158 4048 17174
rect 579613 6626 579679 6629
rect 583520 6626 584960 6716
rect 579613 6624 584960 6626
rect -960 6490 480 6580
rect 579613 6568 579618 6624
rect 579674 6568 584960 6624
rect 579613 6566 584960 6568
rect 579613 6563 579679 6566
rect 2773 6490 2839 6493
rect -960 6488 2839 6490
rect -960 6432 2778 6488
rect 2834 6432 2839 6488
rect 583520 6476 584960 6566
rect -960 6430 2839 6432
rect -960 6340 480 6430
rect 2773 6427 2839 6430
rect 2773 4178 2839 4181
rect 576761 4178 576827 4181
rect 2773 4176 3802 4178
rect 2773 4120 2778 4176
rect 2834 4164 3802 4176
rect 576350 4176 576827 4178
rect 576350 4164 576766 4176
rect 2834 4120 4048 4164
rect 2773 4118 4048 4120
rect 2773 4115 2839 4118
rect 3742 4104 4048 4118
rect 575920 4120 576766 4164
rect 576822 4120 576827 4176
rect 575920 4118 576827 4120
rect 575920 4104 576410 4118
rect 576761 4115 576827 4118
<< metal4 >>
rect -23776 726608 -23156 726640
rect -23776 726372 -23744 726608
rect -23508 726372 -23424 726608
rect -23188 726372 -23156 726608
rect -23776 726288 -23156 726372
rect -23776 726052 -23744 726288
rect -23508 726052 -23424 726288
rect -23188 726052 -23156 726288
rect -23776 669694 -23156 726052
rect -23776 669458 -23744 669694
rect -23508 669458 -23424 669694
rect -23188 669458 -23156 669694
rect -23776 669374 -23156 669458
rect -23776 669138 -23744 669374
rect -23508 669138 -23424 669374
rect -23188 669138 -23156 669374
rect -23776 629694 -23156 669138
rect -23776 629458 -23744 629694
rect -23508 629458 -23424 629694
rect -23188 629458 -23156 629694
rect -23776 629374 -23156 629458
rect -23776 629138 -23744 629374
rect -23508 629138 -23424 629374
rect -23188 629138 -23156 629374
rect -23776 589694 -23156 629138
rect -23776 589458 -23744 589694
rect -23508 589458 -23424 589694
rect -23188 589458 -23156 589694
rect -23776 589374 -23156 589458
rect -23776 589138 -23744 589374
rect -23508 589138 -23424 589374
rect -23188 589138 -23156 589374
rect -23776 549694 -23156 589138
rect -23776 549458 -23744 549694
rect -23508 549458 -23424 549694
rect -23188 549458 -23156 549694
rect -23776 549374 -23156 549458
rect -23776 549138 -23744 549374
rect -23508 549138 -23424 549374
rect -23188 549138 -23156 549374
rect -23776 509694 -23156 549138
rect -23776 509458 -23744 509694
rect -23508 509458 -23424 509694
rect -23188 509458 -23156 509694
rect -23776 509374 -23156 509458
rect -23776 509138 -23744 509374
rect -23508 509138 -23424 509374
rect -23188 509138 -23156 509374
rect -23776 469694 -23156 509138
rect -23776 469458 -23744 469694
rect -23508 469458 -23424 469694
rect -23188 469458 -23156 469694
rect -23776 469374 -23156 469458
rect -23776 469138 -23744 469374
rect -23508 469138 -23424 469374
rect -23188 469138 -23156 469374
rect -23776 429694 -23156 469138
rect -23776 429458 -23744 429694
rect -23508 429458 -23424 429694
rect -23188 429458 -23156 429694
rect -23776 429374 -23156 429458
rect -23776 429138 -23744 429374
rect -23508 429138 -23424 429374
rect -23188 429138 -23156 429374
rect -23776 389694 -23156 429138
rect -23776 389458 -23744 389694
rect -23508 389458 -23424 389694
rect -23188 389458 -23156 389694
rect -23776 389374 -23156 389458
rect -23776 389138 -23744 389374
rect -23508 389138 -23424 389374
rect -23188 389138 -23156 389374
rect -23776 349694 -23156 389138
rect -23776 349458 -23744 349694
rect -23508 349458 -23424 349694
rect -23188 349458 -23156 349694
rect -23776 349374 -23156 349458
rect -23776 349138 -23744 349374
rect -23508 349138 -23424 349374
rect -23188 349138 -23156 349374
rect -23776 309694 -23156 349138
rect -23776 309458 -23744 309694
rect -23508 309458 -23424 309694
rect -23188 309458 -23156 309694
rect -23776 309374 -23156 309458
rect -23776 309138 -23744 309374
rect -23508 309138 -23424 309374
rect -23188 309138 -23156 309374
rect -23776 269694 -23156 309138
rect -23776 269458 -23744 269694
rect -23508 269458 -23424 269694
rect -23188 269458 -23156 269694
rect -23776 269374 -23156 269458
rect -23776 269138 -23744 269374
rect -23508 269138 -23424 269374
rect -23188 269138 -23156 269374
rect -23776 229694 -23156 269138
rect -23776 229458 -23744 229694
rect -23508 229458 -23424 229694
rect -23188 229458 -23156 229694
rect -23776 229374 -23156 229458
rect -23776 229138 -23744 229374
rect -23508 229138 -23424 229374
rect -23188 229138 -23156 229374
rect -23776 189694 -23156 229138
rect -23776 189458 -23744 189694
rect -23508 189458 -23424 189694
rect -23188 189458 -23156 189694
rect -23776 189374 -23156 189458
rect -23776 189138 -23744 189374
rect -23508 189138 -23424 189374
rect -23188 189138 -23156 189374
rect -23776 149694 -23156 189138
rect -23776 149458 -23744 149694
rect -23508 149458 -23424 149694
rect -23188 149458 -23156 149694
rect -23776 149374 -23156 149458
rect -23776 149138 -23744 149374
rect -23508 149138 -23424 149374
rect -23188 149138 -23156 149374
rect -23776 109694 -23156 149138
rect -23776 109458 -23744 109694
rect -23508 109458 -23424 109694
rect -23188 109458 -23156 109694
rect -23776 109374 -23156 109458
rect -23776 109138 -23744 109374
rect -23508 109138 -23424 109374
rect -23188 109138 -23156 109374
rect -23776 69694 -23156 109138
rect -23776 69458 -23744 69694
rect -23508 69458 -23424 69694
rect -23188 69458 -23156 69694
rect -23776 69374 -23156 69458
rect -23776 69138 -23744 69374
rect -23508 69138 -23424 69374
rect -23188 69138 -23156 69374
rect -23776 29694 -23156 69138
rect -23776 29458 -23744 29694
rect -23508 29458 -23424 29694
rect -23188 29458 -23156 29694
rect -23776 29374 -23156 29458
rect -23776 29138 -23744 29374
rect -23508 29138 -23424 29374
rect -23188 29138 -23156 29374
rect -23776 -22116 -23156 29138
rect -20666 723498 -20046 723530
rect -20666 723262 -20634 723498
rect -20398 723262 -20314 723498
rect -20078 723262 -20046 723498
rect -20666 723178 -20046 723262
rect -20666 722942 -20634 723178
rect -20398 722942 -20314 723178
rect -20078 722942 -20046 723178
rect -20666 665974 -20046 722942
rect -20666 665738 -20634 665974
rect -20398 665738 -20314 665974
rect -20078 665738 -20046 665974
rect -20666 665654 -20046 665738
rect -20666 665418 -20634 665654
rect -20398 665418 -20314 665654
rect -20078 665418 -20046 665654
rect -20666 625974 -20046 665418
rect -20666 625738 -20634 625974
rect -20398 625738 -20314 625974
rect -20078 625738 -20046 625974
rect -20666 625654 -20046 625738
rect -20666 625418 -20634 625654
rect -20398 625418 -20314 625654
rect -20078 625418 -20046 625654
rect -20666 585974 -20046 625418
rect -20666 585738 -20634 585974
rect -20398 585738 -20314 585974
rect -20078 585738 -20046 585974
rect -20666 585654 -20046 585738
rect -20666 585418 -20634 585654
rect -20398 585418 -20314 585654
rect -20078 585418 -20046 585654
rect -20666 545974 -20046 585418
rect -20666 545738 -20634 545974
rect -20398 545738 -20314 545974
rect -20078 545738 -20046 545974
rect -20666 545654 -20046 545738
rect -20666 545418 -20634 545654
rect -20398 545418 -20314 545654
rect -20078 545418 -20046 545654
rect -20666 505974 -20046 545418
rect -20666 505738 -20634 505974
rect -20398 505738 -20314 505974
rect -20078 505738 -20046 505974
rect -20666 505654 -20046 505738
rect -20666 505418 -20634 505654
rect -20398 505418 -20314 505654
rect -20078 505418 -20046 505654
rect -20666 465974 -20046 505418
rect -20666 465738 -20634 465974
rect -20398 465738 -20314 465974
rect -20078 465738 -20046 465974
rect -20666 465654 -20046 465738
rect -20666 465418 -20634 465654
rect -20398 465418 -20314 465654
rect -20078 465418 -20046 465654
rect -20666 425974 -20046 465418
rect -20666 425738 -20634 425974
rect -20398 425738 -20314 425974
rect -20078 425738 -20046 425974
rect -20666 425654 -20046 425738
rect -20666 425418 -20634 425654
rect -20398 425418 -20314 425654
rect -20078 425418 -20046 425654
rect -20666 385974 -20046 425418
rect -20666 385738 -20634 385974
rect -20398 385738 -20314 385974
rect -20078 385738 -20046 385974
rect -20666 385654 -20046 385738
rect -20666 385418 -20634 385654
rect -20398 385418 -20314 385654
rect -20078 385418 -20046 385654
rect -20666 345974 -20046 385418
rect -20666 345738 -20634 345974
rect -20398 345738 -20314 345974
rect -20078 345738 -20046 345974
rect -20666 345654 -20046 345738
rect -20666 345418 -20634 345654
rect -20398 345418 -20314 345654
rect -20078 345418 -20046 345654
rect -20666 305974 -20046 345418
rect -20666 305738 -20634 305974
rect -20398 305738 -20314 305974
rect -20078 305738 -20046 305974
rect -20666 305654 -20046 305738
rect -20666 305418 -20634 305654
rect -20398 305418 -20314 305654
rect -20078 305418 -20046 305654
rect -20666 265974 -20046 305418
rect -20666 265738 -20634 265974
rect -20398 265738 -20314 265974
rect -20078 265738 -20046 265974
rect -20666 265654 -20046 265738
rect -20666 265418 -20634 265654
rect -20398 265418 -20314 265654
rect -20078 265418 -20046 265654
rect -20666 225974 -20046 265418
rect -20666 225738 -20634 225974
rect -20398 225738 -20314 225974
rect -20078 225738 -20046 225974
rect -20666 225654 -20046 225738
rect -20666 225418 -20634 225654
rect -20398 225418 -20314 225654
rect -20078 225418 -20046 225654
rect -20666 185974 -20046 225418
rect -20666 185738 -20634 185974
rect -20398 185738 -20314 185974
rect -20078 185738 -20046 185974
rect -20666 185654 -20046 185738
rect -20666 185418 -20634 185654
rect -20398 185418 -20314 185654
rect -20078 185418 -20046 185654
rect -20666 145974 -20046 185418
rect -20666 145738 -20634 145974
rect -20398 145738 -20314 145974
rect -20078 145738 -20046 145974
rect -20666 145654 -20046 145738
rect -20666 145418 -20634 145654
rect -20398 145418 -20314 145654
rect -20078 145418 -20046 145654
rect -20666 105974 -20046 145418
rect -20666 105738 -20634 105974
rect -20398 105738 -20314 105974
rect -20078 105738 -20046 105974
rect -20666 105654 -20046 105738
rect -20666 105418 -20634 105654
rect -20398 105418 -20314 105654
rect -20078 105418 -20046 105654
rect -20666 65974 -20046 105418
rect -20666 65738 -20634 65974
rect -20398 65738 -20314 65974
rect -20078 65738 -20046 65974
rect -20666 65654 -20046 65738
rect -20666 65418 -20634 65654
rect -20398 65418 -20314 65654
rect -20078 65418 -20046 65654
rect -20666 25974 -20046 65418
rect -20666 25738 -20634 25974
rect -20398 25738 -20314 25974
rect -20078 25738 -20046 25974
rect -20666 25654 -20046 25738
rect -20666 25418 -20634 25654
rect -20398 25418 -20314 25654
rect -20078 25418 -20046 25654
rect -20666 -19006 -20046 25418
rect -17556 720388 -16936 720420
rect -17556 720152 -17524 720388
rect -17288 720152 -17204 720388
rect -16968 720152 -16936 720388
rect -17556 720068 -16936 720152
rect -17556 719832 -17524 720068
rect -17288 719832 -17204 720068
rect -16968 719832 -16936 720068
rect -17556 662254 -16936 719832
rect 580594 720388 581214 726640
rect 607080 726608 607700 726640
rect 607080 726372 607112 726608
rect 607348 726372 607432 726608
rect 607668 726372 607700 726608
rect 607080 726288 607700 726372
rect 607080 726052 607112 726288
rect 607348 726052 607432 726288
rect 607668 726052 607700 726288
rect 603970 723498 604590 723530
rect 603970 723262 604002 723498
rect 604238 723262 604322 723498
rect 604558 723262 604590 723498
rect 603970 723178 604590 723262
rect 603970 722942 604002 723178
rect 604238 722942 604322 723178
rect 604558 722942 604590 723178
rect 580594 720152 580626 720388
rect 580862 720152 580946 720388
rect 581182 720152 581214 720388
rect 580594 720068 581214 720152
rect 580594 719832 580626 720068
rect 580862 719832 580946 720068
rect 581182 719832 581214 720068
rect -17556 662018 -17524 662254
rect -17288 662018 -17204 662254
rect -16968 662018 -16936 662254
rect -17556 661934 -16936 662018
rect -17556 661698 -17524 661934
rect -17288 661698 -17204 661934
rect -16968 661698 -16936 661934
rect -17556 622254 -16936 661698
rect -17556 622018 -17524 622254
rect -17288 622018 -17204 622254
rect -16968 622018 -16936 622254
rect -17556 621934 -16936 622018
rect -17556 621698 -17524 621934
rect -17288 621698 -17204 621934
rect -16968 621698 -16936 621934
rect -17556 582254 -16936 621698
rect -17556 582018 -17524 582254
rect -17288 582018 -17204 582254
rect -16968 582018 -16936 582254
rect -17556 581934 -16936 582018
rect -17556 581698 -17524 581934
rect -17288 581698 -17204 581934
rect -16968 581698 -16936 581934
rect -17556 542254 -16936 581698
rect -17556 542018 -17524 542254
rect -17288 542018 -17204 542254
rect -16968 542018 -16936 542254
rect -17556 541934 -16936 542018
rect -17556 541698 -17524 541934
rect -17288 541698 -17204 541934
rect -16968 541698 -16936 541934
rect -17556 502254 -16936 541698
rect -17556 502018 -17524 502254
rect -17288 502018 -17204 502254
rect -16968 502018 -16936 502254
rect -17556 501934 -16936 502018
rect -17556 501698 -17524 501934
rect -17288 501698 -17204 501934
rect -16968 501698 -16936 501934
rect -17556 462254 -16936 501698
rect -17556 462018 -17524 462254
rect -17288 462018 -17204 462254
rect -16968 462018 -16936 462254
rect -17556 461934 -16936 462018
rect -17556 461698 -17524 461934
rect -17288 461698 -17204 461934
rect -16968 461698 -16936 461934
rect -17556 422254 -16936 461698
rect -17556 422018 -17524 422254
rect -17288 422018 -17204 422254
rect -16968 422018 -16936 422254
rect -17556 421934 -16936 422018
rect -17556 421698 -17524 421934
rect -17288 421698 -17204 421934
rect -16968 421698 -16936 421934
rect -17556 382254 -16936 421698
rect -17556 382018 -17524 382254
rect -17288 382018 -17204 382254
rect -16968 382018 -16936 382254
rect -17556 381934 -16936 382018
rect -17556 381698 -17524 381934
rect -17288 381698 -17204 381934
rect -16968 381698 -16936 381934
rect -17556 342254 -16936 381698
rect -17556 342018 -17524 342254
rect -17288 342018 -17204 342254
rect -16968 342018 -16936 342254
rect -17556 341934 -16936 342018
rect -17556 341698 -17524 341934
rect -17288 341698 -17204 341934
rect -16968 341698 -16936 341934
rect -17556 302254 -16936 341698
rect -17556 302018 -17524 302254
rect -17288 302018 -17204 302254
rect -16968 302018 -16936 302254
rect -17556 301934 -16936 302018
rect -17556 301698 -17524 301934
rect -17288 301698 -17204 301934
rect -16968 301698 -16936 301934
rect -17556 262254 -16936 301698
rect -17556 262018 -17524 262254
rect -17288 262018 -17204 262254
rect -16968 262018 -16936 262254
rect -17556 261934 -16936 262018
rect -17556 261698 -17524 261934
rect -17288 261698 -17204 261934
rect -16968 261698 -16936 261934
rect -17556 222254 -16936 261698
rect -17556 222018 -17524 222254
rect -17288 222018 -17204 222254
rect -16968 222018 -16936 222254
rect -17556 221934 -16936 222018
rect -17556 221698 -17524 221934
rect -17288 221698 -17204 221934
rect -16968 221698 -16936 221934
rect -17556 182254 -16936 221698
rect -17556 182018 -17524 182254
rect -17288 182018 -17204 182254
rect -16968 182018 -16936 182254
rect -17556 181934 -16936 182018
rect -17556 181698 -17524 181934
rect -17288 181698 -17204 181934
rect -16968 181698 -16936 181934
rect -17556 142254 -16936 181698
rect -17556 142018 -17524 142254
rect -17288 142018 -17204 142254
rect -16968 142018 -16936 142254
rect -17556 141934 -16936 142018
rect -17556 141698 -17524 141934
rect -17288 141698 -17204 141934
rect -16968 141698 -16936 141934
rect -17556 102254 -16936 141698
rect -17556 102018 -17524 102254
rect -17288 102018 -17204 102254
rect -16968 102018 -16936 102254
rect -17556 101934 -16936 102018
rect -17556 101698 -17524 101934
rect -17288 101698 -17204 101934
rect -16968 101698 -16936 101934
rect -17556 62254 -16936 101698
rect -17556 62018 -17524 62254
rect -17288 62018 -17204 62254
rect -16968 62018 -16936 62254
rect -17556 61934 -16936 62018
rect -17556 61698 -17524 61934
rect -17288 61698 -17204 61934
rect -16968 61698 -16936 61934
rect -17556 22254 -16936 61698
rect -17556 22018 -17524 22254
rect -17288 22018 -17204 22254
rect -16968 22018 -16936 22254
rect -17556 21934 -16936 22018
rect -17556 21698 -17524 21934
rect -17288 21698 -17204 21934
rect -16968 21698 -16936 21934
rect -17556 -15896 -16936 21698
rect -14446 717278 -13826 717310
rect -14446 717042 -14414 717278
rect -14178 717042 -14094 717278
rect -13858 717042 -13826 717278
rect -14446 716958 -13826 717042
rect -14446 716722 -14414 716958
rect -14178 716722 -14094 716958
rect -13858 716722 -13826 716958
rect -14446 698534 -13826 716722
rect -14446 698298 -14414 698534
rect -14178 698298 -14094 698534
rect -13858 698298 -13826 698534
rect -14446 698214 -13826 698298
rect -14446 697978 -14414 698214
rect -14178 697978 -14094 698214
rect -13858 697978 -13826 698214
rect -14446 658534 -13826 697978
rect -14446 658298 -14414 658534
rect -14178 658298 -14094 658534
rect -13858 658298 -13826 658534
rect -14446 658214 -13826 658298
rect -14446 657978 -14414 658214
rect -14178 657978 -14094 658214
rect -13858 657978 -13826 658214
rect -14446 618534 -13826 657978
rect -14446 618298 -14414 618534
rect -14178 618298 -14094 618534
rect -13858 618298 -13826 618534
rect -14446 618214 -13826 618298
rect -14446 617978 -14414 618214
rect -14178 617978 -14094 618214
rect -13858 617978 -13826 618214
rect -14446 578534 -13826 617978
rect -14446 578298 -14414 578534
rect -14178 578298 -14094 578534
rect -13858 578298 -13826 578534
rect -14446 578214 -13826 578298
rect -14446 577978 -14414 578214
rect -14178 577978 -14094 578214
rect -13858 577978 -13826 578214
rect -14446 538534 -13826 577978
rect -14446 538298 -14414 538534
rect -14178 538298 -14094 538534
rect -13858 538298 -13826 538534
rect -14446 538214 -13826 538298
rect -14446 537978 -14414 538214
rect -14178 537978 -14094 538214
rect -13858 537978 -13826 538214
rect -14446 498534 -13826 537978
rect -14446 498298 -14414 498534
rect -14178 498298 -14094 498534
rect -13858 498298 -13826 498534
rect -14446 498214 -13826 498298
rect -14446 497978 -14414 498214
rect -14178 497978 -14094 498214
rect -13858 497978 -13826 498214
rect -14446 458534 -13826 497978
rect -14446 458298 -14414 458534
rect -14178 458298 -14094 458534
rect -13858 458298 -13826 458534
rect -14446 458214 -13826 458298
rect -14446 457978 -14414 458214
rect -14178 457978 -14094 458214
rect -13858 457978 -13826 458214
rect -14446 418534 -13826 457978
rect -14446 418298 -14414 418534
rect -14178 418298 -14094 418534
rect -13858 418298 -13826 418534
rect -14446 418214 -13826 418298
rect -14446 417978 -14414 418214
rect -14178 417978 -14094 418214
rect -13858 417978 -13826 418214
rect -14446 378534 -13826 417978
rect -14446 378298 -14414 378534
rect -14178 378298 -14094 378534
rect -13858 378298 -13826 378534
rect -14446 378214 -13826 378298
rect -14446 377978 -14414 378214
rect -14178 377978 -14094 378214
rect -13858 377978 -13826 378214
rect -14446 338534 -13826 377978
rect -14446 338298 -14414 338534
rect -14178 338298 -14094 338534
rect -13858 338298 -13826 338534
rect -14446 338214 -13826 338298
rect -14446 337978 -14414 338214
rect -14178 337978 -14094 338214
rect -13858 337978 -13826 338214
rect -14446 298534 -13826 337978
rect -14446 298298 -14414 298534
rect -14178 298298 -14094 298534
rect -13858 298298 -13826 298534
rect -14446 298214 -13826 298298
rect -14446 297978 -14414 298214
rect -14178 297978 -14094 298214
rect -13858 297978 -13826 298214
rect -14446 258534 -13826 297978
rect -14446 258298 -14414 258534
rect -14178 258298 -14094 258534
rect -13858 258298 -13826 258534
rect -14446 258214 -13826 258298
rect -14446 257978 -14414 258214
rect -14178 257978 -14094 258214
rect -13858 257978 -13826 258214
rect -14446 218534 -13826 257978
rect -14446 218298 -14414 218534
rect -14178 218298 -14094 218534
rect -13858 218298 -13826 218534
rect -14446 218214 -13826 218298
rect -14446 217978 -14414 218214
rect -14178 217978 -14094 218214
rect -13858 217978 -13826 218214
rect -14446 178534 -13826 217978
rect -14446 178298 -14414 178534
rect -14178 178298 -14094 178534
rect -13858 178298 -13826 178534
rect -14446 178214 -13826 178298
rect -14446 177978 -14414 178214
rect -14178 177978 -14094 178214
rect -13858 177978 -13826 178214
rect -14446 138534 -13826 177978
rect -14446 138298 -14414 138534
rect -14178 138298 -14094 138534
rect -13858 138298 -13826 138534
rect -14446 138214 -13826 138298
rect -14446 137978 -14414 138214
rect -14178 137978 -14094 138214
rect -13858 137978 -13826 138214
rect -14446 98534 -13826 137978
rect -14446 98298 -14414 98534
rect -14178 98298 -14094 98534
rect -13858 98298 -13826 98534
rect -14446 98214 -13826 98298
rect -14446 97978 -14414 98214
rect -14178 97978 -14094 98214
rect -13858 97978 -13826 98214
rect -14446 58534 -13826 97978
rect -14446 58298 -14414 58534
rect -14178 58298 -14094 58534
rect -13858 58298 -13826 58534
rect -14446 58214 -13826 58298
rect -14446 57978 -14414 58214
rect -14178 57978 -14094 58214
rect -13858 57978 -13826 58214
rect -14446 18534 -13826 57978
rect -14446 18298 -14414 18534
rect -14178 18298 -14094 18534
rect -13858 18298 -13826 18534
rect -14446 18214 -13826 18298
rect -14446 17978 -14414 18214
rect -14178 17978 -14094 18214
rect -13858 17978 -13826 18214
rect -14446 -12786 -13826 17978
rect -11336 714168 -10716 714200
rect -11336 713932 -11304 714168
rect -11068 713932 -10984 714168
rect -10748 713932 -10716 714168
rect -11336 713848 -10716 713932
rect -11336 713612 -11304 713848
rect -11068 713612 -10984 713848
rect -10748 713612 -10716 713848
rect -11336 694814 -10716 713612
rect -11336 694578 -11304 694814
rect -11068 694578 -10984 694814
rect -10748 694578 -10716 694814
rect -11336 694494 -10716 694578
rect -11336 694258 -11304 694494
rect -11068 694258 -10984 694494
rect -10748 694258 -10716 694494
rect -11336 654814 -10716 694258
rect -11336 654578 -11304 654814
rect -11068 654578 -10984 654814
rect -10748 654578 -10716 654814
rect -11336 654494 -10716 654578
rect -11336 654258 -11304 654494
rect -11068 654258 -10984 654494
rect -10748 654258 -10716 654494
rect -11336 614814 -10716 654258
rect -11336 614578 -11304 614814
rect -11068 614578 -10984 614814
rect -10748 614578 -10716 614814
rect -11336 614494 -10716 614578
rect -11336 614258 -11304 614494
rect -11068 614258 -10984 614494
rect -10748 614258 -10716 614494
rect -11336 574814 -10716 614258
rect -11336 574578 -11304 574814
rect -11068 574578 -10984 574814
rect -10748 574578 -10716 574814
rect -11336 574494 -10716 574578
rect -11336 574258 -11304 574494
rect -11068 574258 -10984 574494
rect -10748 574258 -10716 574494
rect -11336 534814 -10716 574258
rect -11336 534578 -11304 534814
rect -11068 534578 -10984 534814
rect -10748 534578 -10716 534814
rect -11336 534494 -10716 534578
rect -11336 534258 -11304 534494
rect -11068 534258 -10984 534494
rect -10748 534258 -10716 534494
rect -11336 494814 -10716 534258
rect -11336 494578 -11304 494814
rect -11068 494578 -10984 494814
rect -10748 494578 -10716 494814
rect -11336 494494 -10716 494578
rect -11336 494258 -11304 494494
rect -11068 494258 -10984 494494
rect -10748 494258 -10716 494494
rect -11336 454814 -10716 494258
rect -11336 454578 -11304 454814
rect -11068 454578 -10984 454814
rect -10748 454578 -10716 454814
rect -11336 454494 -10716 454578
rect -11336 454258 -11304 454494
rect -11068 454258 -10984 454494
rect -10748 454258 -10716 454494
rect -11336 414814 -10716 454258
rect -11336 414578 -11304 414814
rect -11068 414578 -10984 414814
rect -10748 414578 -10716 414814
rect -11336 414494 -10716 414578
rect -11336 414258 -11304 414494
rect -11068 414258 -10984 414494
rect -10748 414258 -10716 414494
rect -11336 374814 -10716 414258
rect -11336 374578 -11304 374814
rect -11068 374578 -10984 374814
rect -10748 374578 -10716 374814
rect -11336 374494 -10716 374578
rect -11336 374258 -11304 374494
rect -11068 374258 -10984 374494
rect -10748 374258 -10716 374494
rect -11336 334814 -10716 374258
rect -11336 334578 -11304 334814
rect -11068 334578 -10984 334814
rect -10748 334578 -10716 334814
rect -11336 334494 -10716 334578
rect -11336 334258 -11304 334494
rect -11068 334258 -10984 334494
rect -10748 334258 -10716 334494
rect -11336 294814 -10716 334258
rect -11336 294578 -11304 294814
rect -11068 294578 -10984 294814
rect -10748 294578 -10716 294814
rect -11336 294494 -10716 294578
rect -11336 294258 -11304 294494
rect -11068 294258 -10984 294494
rect -10748 294258 -10716 294494
rect -11336 254814 -10716 294258
rect -11336 254578 -11304 254814
rect -11068 254578 -10984 254814
rect -10748 254578 -10716 254814
rect -11336 254494 -10716 254578
rect -11336 254258 -11304 254494
rect -11068 254258 -10984 254494
rect -10748 254258 -10716 254494
rect -11336 214814 -10716 254258
rect -11336 214578 -11304 214814
rect -11068 214578 -10984 214814
rect -10748 214578 -10716 214814
rect -11336 214494 -10716 214578
rect -11336 214258 -11304 214494
rect -11068 214258 -10984 214494
rect -10748 214258 -10716 214494
rect -11336 174814 -10716 214258
rect -11336 174578 -11304 174814
rect -11068 174578 -10984 174814
rect -10748 174578 -10716 174814
rect -11336 174494 -10716 174578
rect -11336 174258 -11304 174494
rect -11068 174258 -10984 174494
rect -10748 174258 -10716 174494
rect -11336 134814 -10716 174258
rect -11336 134578 -11304 134814
rect -11068 134578 -10984 134814
rect -10748 134578 -10716 134814
rect -11336 134494 -10716 134578
rect -11336 134258 -11304 134494
rect -11068 134258 -10984 134494
rect -10748 134258 -10716 134494
rect -11336 94814 -10716 134258
rect -11336 94578 -11304 94814
rect -11068 94578 -10984 94814
rect -10748 94578 -10716 94814
rect -11336 94494 -10716 94578
rect -11336 94258 -11304 94494
rect -11068 94258 -10984 94494
rect -10748 94258 -10716 94494
rect -11336 54814 -10716 94258
rect -11336 54578 -11304 54814
rect -11068 54578 -10984 54814
rect -10748 54578 -10716 54814
rect -11336 54494 -10716 54578
rect -11336 54258 -11304 54494
rect -11068 54258 -10984 54494
rect -10748 54258 -10716 54494
rect -11336 14814 -10716 54258
rect -11336 14578 -11304 14814
rect -11068 14578 -10984 14814
rect -10748 14578 -10716 14814
rect -11336 14494 -10716 14578
rect -11336 14258 -11304 14494
rect -11068 14258 -10984 14494
rect -10748 14258 -10716 14494
rect -11336 -9676 -10716 14258
rect -8226 711058 -7606 711090
rect -8226 710822 -8194 711058
rect -7958 710822 -7874 711058
rect -7638 710822 -7606 711058
rect -8226 710738 -7606 710822
rect -8226 710502 -8194 710738
rect -7958 710502 -7874 710738
rect -7638 710502 -7606 710738
rect -8226 691094 -7606 710502
rect -8226 690858 -8194 691094
rect -7958 690858 -7874 691094
rect -7638 690858 -7606 691094
rect -8226 690774 -7606 690858
rect -8226 690538 -8194 690774
rect -7958 690538 -7874 690774
rect -7638 690538 -7606 690774
rect -8226 651094 -7606 690538
rect -8226 650858 -8194 651094
rect -7958 650858 -7874 651094
rect -7638 650858 -7606 651094
rect -8226 650774 -7606 650858
rect -8226 650538 -8194 650774
rect -7958 650538 -7874 650774
rect -7638 650538 -7606 650774
rect -8226 611094 -7606 650538
rect -8226 610858 -8194 611094
rect -7958 610858 -7874 611094
rect -7638 610858 -7606 611094
rect -8226 610774 -7606 610858
rect -8226 610538 -8194 610774
rect -7958 610538 -7874 610774
rect -7638 610538 -7606 610774
rect -8226 571094 -7606 610538
rect -8226 570858 -8194 571094
rect -7958 570858 -7874 571094
rect -7638 570858 -7606 571094
rect -8226 570774 -7606 570858
rect -8226 570538 -8194 570774
rect -7958 570538 -7874 570774
rect -7638 570538 -7606 570774
rect -8226 531094 -7606 570538
rect -8226 530858 -8194 531094
rect -7958 530858 -7874 531094
rect -7638 530858 -7606 531094
rect -8226 530774 -7606 530858
rect -8226 530538 -8194 530774
rect -7958 530538 -7874 530774
rect -7638 530538 -7606 530774
rect -8226 491094 -7606 530538
rect -8226 490858 -8194 491094
rect -7958 490858 -7874 491094
rect -7638 490858 -7606 491094
rect -8226 490774 -7606 490858
rect -8226 490538 -8194 490774
rect -7958 490538 -7874 490774
rect -7638 490538 -7606 490774
rect -8226 451094 -7606 490538
rect -8226 450858 -8194 451094
rect -7958 450858 -7874 451094
rect -7638 450858 -7606 451094
rect -8226 450774 -7606 450858
rect -8226 450538 -8194 450774
rect -7958 450538 -7874 450774
rect -7638 450538 -7606 450774
rect -8226 411094 -7606 450538
rect -8226 410858 -8194 411094
rect -7958 410858 -7874 411094
rect -7638 410858 -7606 411094
rect -8226 410774 -7606 410858
rect -8226 410538 -8194 410774
rect -7958 410538 -7874 410774
rect -7638 410538 -7606 410774
rect -8226 371094 -7606 410538
rect -8226 370858 -8194 371094
rect -7958 370858 -7874 371094
rect -7638 370858 -7606 371094
rect -8226 370774 -7606 370858
rect -8226 370538 -8194 370774
rect -7958 370538 -7874 370774
rect -7638 370538 -7606 370774
rect -8226 331094 -7606 370538
rect -8226 330858 -8194 331094
rect -7958 330858 -7874 331094
rect -7638 330858 -7606 331094
rect -8226 330774 -7606 330858
rect -8226 330538 -8194 330774
rect -7958 330538 -7874 330774
rect -7638 330538 -7606 330774
rect -8226 291094 -7606 330538
rect -8226 290858 -8194 291094
rect -7958 290858 -7874 291094
rect -7638 290858 -7606 291094
rect -8226 290774 -7606 290858
rect -8226 290538 -8194 290774
rect -7958 290538 -7874 290774
rect -7638 290538 -7606 290774
rect -8226 251094 -7606 290538
rect -8226 250858 -8194 251094
rect -7958 250858 -7874 251094
rect -7638 250858 -7606 251094
rect -8226 250774 -7606 250858
rect -8226 250538 -8194 250774
rect -7958 250538 -7874 250774
rect -7638 250538 -7606 250774
rect -8226 211094 -7606 250538
rect -8226 210858 -8194 211094
rect -7958 210858 -7874 211094
rect -7638 210858 -7606 211094
rect -8226 210774 -7606 210858
rect -8226 210538 -8194 210774
rect -7958 210538 -7874 210774
rect -7638 210538 -7606 210774
rect -8226 171094 -7606 210538
rect -8226 170858 -8194 171094
rect -7958 170858 -7874 171094
rect -7638 170858 -7606 171094
rect -8226 170774 -7606 170858
rect -8226 170538 -8194 170774
rect -7958 170538 -7874 170774
rect -7638 170538 -7606 170774
rect -8226 131094 -7606 170538
rect -8226 130858 -8194 131094
rect -7958 130858 -7874 131094
rect -7638 130858 -7606 131094
rect -8226 130774 -7606 130858
rect -8226 130538 -8194 130774
rect -7958 130538 -7874 130774
rect -7638 130538 -7606 130774
rect -8226 91094 -7606 130538
rect -8226 90858 -8194 91094
rect -7958 90858 -7874 91094
rect -7638 90858 -7606 91094
rect -8226 90774 -7606 90858
rect -8226 90538 -8194 90774
rect -7958 90538 -7874 90774
rect -7638 90538 -7606 90774
rect -8226 51094 -7606 90538
rect -8226 50858 -8194 51094
rect -7958 50858 -7874 51094
rect -7638 50858 -7606 51094
rect -8226 50774 -7606 50858
rect -8226 50538 -8194 50774
rect -7958 50538 -7874 50774
rect -7638 50538 -7606 50774
rect -8226 11094 -7606 50538
rect -8226 10858 -8194 11094
rect -7958 10858 -7874 11094
rect -7638 10858 -7606 11094
rect -8226 10774 -7606 10858
rect -8226 10538 -8194 10774
rect -7958 10538 -7874 10774
rect -7638 10538 -7606 10774
rect -8226 -6566 -7606 10538
rect -5116 707948 -4496 707980
rect -5116 707712 -5084 707948
rect -4848 707712 -4764 707948
rect -4528 707712 -4496 707948
rect -5116 707628 -4496 707712
rect -5116 707392 -5084 707628
rect -4848 707392 -4764 707628
rect -4528 707392 -4496 707628
rect -5116 687374 -4496 707392
rect -5116 687138 -5084 687374
rect -4848 687138 -4764 687374
rect -4528 687138 -4496 687374
rect -5116 687054 -4496 687138
rect -5116 686818 -5084 687054
rect -4848 686818 -4764 687054
rect -4528 686818 -4496 687054
rect -5116 647374 -4496 686818
rect -5116 647138 -5084 647374
rect -4848 647138 -4764 647374
rect -4528 647138 -4496 647374
rect -5116 647054 -4496 647138
rect -5116 646818 -5084 647054
rect -4848 646818 -4764 647054
rect -4528 646818 -4496 647054
rect -5116 607374 -4496 646818
rect -5116 607138 -5084 607374
rect -4848 607138 -4764 607374
rect -4528 607138 -4496 607374
rect -5116 607054 -4496 607138
rect -5116 606818 -5084 607054
rect -4848 606818 -4764 607054
rect -4528 606818 -4496 607054
rect -5116 567374 -4496 606818
rect -5116 567138 -5084 567374
rect -4848 567138 -4764 567374
rect -4528 567138 -4496 567374
rect -5116 567054 -4496 567138
rect -5116 566818 -5084 567054
rect -4848 566818 -4764 567054
rect -4528 566818 -4496 567054
rect -5116 527374 -4496 566818
rect -5116 527138 -5084 527374
rect -4848 527138 -4764 527374
rect -4528 527138 -4496 527374
rect -5116 527054 -4496 527138
rect -5116 526818 -5084 527054
rect -4848 526818 -4764 527054
rect -4528 526818 -4496 527054
rect -5116 487374 -4496 526818
rect -5116 487138 -5084 487374
rect -4848 487138 -4764 487374
rect -4528 487138 -4496 487374
rect -5116 487054 -4496 487138
rect -5116 486818 -5084 487054
rect -4848 486818 -4764 487054
rect -4528 486818 -4496 487054
rect -5116 447374 -4496 486818
rect -5116 447138 -5084 447374
rect -4848 447138 -4764 447374
rect -4528 447138 -4496 447374
rect -5116 447054 -4496 447138
rect -5116 446818 -5084 447054
rect -4848 446818 -4764 447054
rect -4528 446818 -4496 447054
rect -5116 407374 -4496 446818
rect -5116 407138 -5084 407374
rect -4848 407138 -4764 407374
rect -4528 407138 -4496 407374
rect -5116 407054 -4496 407138
rect -5116 406818 -5084 407054
rect -4848 406818 -4764 407054
rect -4528 406818 -4496 407054
rect -5116 367374 -4496 406818
rect -5116 367138 -5084 367374
rect -4848 367138 -4764 367374
rect -4528 367138 -4496 367374
rect -5116 367054 -4496 367138
rect -5116 366818 -5084 367054
rect -4848 366818 -4764 367054
rect -4528 366818 -4496 367054
rect -5116 327374 -4496 366818
rect -5116 327138 -5084 327374
rect -4848 327138 -4764 327374
rect -4528 327138 -4496 327374
rect -5116 327054 -4496 327138
rect -5116 326818 -5084 327054
rect -4848 326818 -4764 327054
rect -4528 326818 -4496 327054
rect -5116 287374 -4496 326818
rect -5116 287138 -5084 287374
rect -4848 287138 -4764 287374
rect -4528 287138 -4496 287374
rect -5116 287054 -4496 287138
rect -5116 286818 -5084 287054
rect -4848 286818 -4764 287054
rect -4528 286818 -4496 287054
rect -5116 247374 -4496 286818
rect -5116 247138 -5084 247374
rect -4848 247138 -4764 247374
rect -4528 247138 -4496 247374
rect -5116 247054 -4496 247138
rect -5116 246818 -5084 247054
rect -4848 246818 -4764 247054
rect -4528 246818 -4496 247054
rect -5116 207374 -4496 246818
rect -5116 207138 -5084 207374
rect -4848 207138 -4764 207374
rect -4528 207138 -4496 207374
rect -5116 207054 -4496 207138
rect -5116 206818 -5084 207054
rect -4848 206818 -4764 207054
rect -4528 206818 -4496 207054
rect -5116 167374 -4496 206818
rect -5116 167138 -5084 167374
rect -4848 167138 -4764 167374
rect -4528 167138 -4496 167374
rect -5116 167054 -4496 167138
rect -5116 166818 -5084 167054
rect -4848 166818 -4764 167054
rect -4528 166818 -4496 167054
rect -5116 127374 -4496 166818
rect -5116 127138 -5084 127374
rect -4848 127138 -4764 127374
rect -4528 127138 -4496 127374
rect -5116 127054 -4496 127138
rect -5116 126818 -5084 127054
rect -4848 126818 -4764 127054
rect -4528 126818 -4496 127054
rect -5116 87374 -4496 126818
rect -5116 87138 -5084 87374
rect -4848 87138 -4764 87374
rect -4528 87138 -4496 87374
rect -5116 87054 -4496 87138
rect -5116 86818 -5084 87054
rect -4848 86818 -4764 87054
rect -4528 86818 -4496 87054
rect -5116 47374 -4496 86818
rect -5116 47138 -5084 47374
rect -4848 47138 -4764 47374
rect -4528 47138 -4496 47374
rect -5116 47054 -4496 47138
rect -5116 46818 -5084 47054
rect -4848 46818 -4764 47054
rect -4528 46818 -4496 47054
rect -5116 7374 -4496 46818
rect -5116 7138 -5084 7374
rect -4848 7138 -4764 7374
rect -4528 7138 -4496 7374
rect -5116 7054 -4496 7138
rect -5116 6818 -5084 7054
rect -4848 6818 -4764 7054
rect -4528 6818 -4496 7054
rect -5116 -3456 -4496 6818
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 683654 -1386 704282
rect 7844 693480 7876 693716
rect 8112 693480 8196 693716
rect 8432 693480 8464 693716
rect 7844 693396 8464 693480
rect 7844 693160 7876 693396
rect 8112 693160 8196 693396
rect 8432 693160 8464 693396
rect 38000 693480 38032 693716
rect 38268 693480 38352 693716
rect 38588 693480 38620 693716
rect 38000 693396 38620 693480
rect 38000 693160 38032 693396
rect 38268 693160 38352 693396
rect 38588 693160 38620 693396
rect 74000 693480 74032 693716
rect 74268 693480 74352 693716
rect 74588 693480 74620 693716
rect 74000 693396 74620 693480
rect 74000 693160 74032 693396
rect 74268 693160 74352 693396
rect 74588 693160 74620 693396
rect 110000 693480 110032 693716
rect 110268 693480 110352 693716
rect 110588 693480 110620 693716
rect 110000 693396 110620 693480
rect 110000 693160 110032 693396
rect 110268 693160 110352 693396
rect 110588 693160 110620 693396
rect 146000 693480 146032 693716
rect 146268 693480 146352 693716
rect 146588 693480 146620 693716
rect 146000 693396 146620 693480
rect 146000 693160 146032 693396
rect 146268 693160 146352 693396
rect 146588 693160 146620 693396
rect 182000 693480 182032 693716
rect 182268 693480 182352 693716
rect 182588 693480 182620 693716
rect 182000 693396 182620 693480
rect 182000 693160 182032 693396
rect 182268 693160 182352 693396
rect 182588 693160 182620 693396
rect 218000 693480 218032 693716
rect 218268 693480 218352 693716
rect 218588 693480 218620 693716
rect 218000 693396 218620 693480
rect 218000 693160 218032 693396
rect 218268 693160 218352 693396
rect 218588 693160 218620 693396
rect 254000 693480 254032 693716
rect 254268 693480 254352 693716
rect 254588 693480 254620 693716
rect 254000 693396 254620 693480
rect 254000 693160 254032 693396
rect 254268 693160 254352 693396
rect 254588 693160 254620 693396
rect 290000 693480 290032 693716
rect 290268 693480 290352 693716
rect 290588 693480 290620 693716
rect 290000 693396 290620 693480
rect 290000 693160 290032 693396
rect 290268 693160 290352 693396
rect 290588 693160 290620 693396
rect 326000 693480 326032 693716
rect 326268 693480 326352 693716
rect 326588 693480 326620 693716
rect 326000 693396 326620 693480
rect 326000 693160 326032 693396
rect 326268 693160 326352 693396
rect 326588 693160 326620 693396
rect 362000 693480 362032 693716
rect 362268 693480 362352 693716
rect 362588 693480 362620 693716
rect 362000 693396 362620 693480
rect 362000 693160 362032 693396
rect 362268 693160 362352 693396
rect 362588 693160 362620 693396
rect 398000 693480 398032 693716
rect 398268 693480 398352 693716
rect 398588 693480 398620 693716
rect 398000 693396 398620 693480
rect 398000 693160 398032 693396
rect 398268 693160 398352 693396
rect 398588 693160 398620 693396
rect 434000 693480 434032 693716
rect 434268 693480 434352 693716
rect 434588 693480 434620 693716
rect 434000 693396 434620 693480
rect 434000 693160 434032 693396
rect 434268 693160 434352 693396
rect 434588 693160 434620 693396
rect 470000 693480 470032 693716
rect 470268 693480 470352 693716
rect 470588 693480 470620 693716
rect 470000 693396 470620 693480
rect 470000 693160 470032 693396
rect 470268 693160 470352 693396
rect 470588 693160 470620 693396
rect 506000 693480 506032 693716
rect 506268 693480 506352 693716
rect 506588 693480 506620 693716
rect 506000 693396 506620 693480
rect 506000 693160 506032 693396
rect 506268 693160 506352 693396
rect 506588 693160 506620 693396
rect 542000 693480 542032 693716
rect 542268 693480 542352 693716
rect 542588 693480 542620 693716
rect 542000 693396 542620 693480
rect 542000 693160 542032 693396
rect 542268 693160 542352 693396
rect 542588 693160 542620 693396
rect 571500 693480 571532 693716
rect 571768 693480 571852 693716
rect 572088 693480 572120 693716
rect 571500 693396 572120 693480
rect 571500 693160 571532 693396
rect 571768 693160 571852 693396
rect 572088 693160 572120 693396
rect 9084 692240 9116 692476
rect 9352 692240 9436 692476
rect 9672 692240 9704 692476
rect 9084 692156 9704 692240
rect 9084 691920 9116 692156
rect 9352 691920 9436 692156
rect 9672 691920 9704 692156
rect 56620 692240 56652 692476
rect 56888 692240 56972 692476
rect 57208 692240 57240 692476
rect 56620 692156 57240 692240
rect 56620 691920 56652 692156
rect 56888 691920 56972 692156
rect 57208 691920 57240 692156
rect 92620 692240 92652 692476
rect 92888 692240 92972 692476
rect 93208 692240 93240 692476
rect 92620 692156 93240 692240
rect 92620 691920 92652 692156
rect 92888 691920 92972 692156
rect 93208 691920 93240 692156
rect 128620 692240 128652 692476
rect 128888 692240 128972 692476
rect 129208 692240 129240 692476
rect 128620 692156 129240 692240
rect 128620 691920 128652 692156
rect 128888 691920 128972 692156
rect 129208 691920 129240 692156
rect 164620 692240 164652 692476
rect 164888 692240 164972 692476
rect 165208 692240 165240 692476
rect 164620 692156 165240 692240
rect 164620 691920 164652 692156
rect 164888 691920 164972 692156
rect 165208 691920 165240 692156
rect 200620 692240 200652 692476
rect 200888 692240 200972 692476
rect 201208 692240 201240 692476
rect 200620 692156 201240 692240
rect 200620 691920 200652 692156
rect 200888 691920 200972 692156
rect 201208 691920 201240 692156
rect 236620 692240 236652 692476
rect 236888 692240 236972 692476
rect 237208 692240 237240 692476
rect 236620 692156 237240 692240
rect 236620 691920 236652 692156
rect 236888 691920 236972 692156
rect 237208 691920 237240 692156
rect 272620 692240 272652 692476
rect 272888 692240 272972 692476
rect 273208 692240 273240 692476
rect 272620 692156 273240 692240
rect 272620 691920 272652 692156
rect 272888 691920 272972 692156
rect 273208 691920 273240 692156
rect 308620 692240 308652 692476
rect 308888 692240 308972 692476
rect 309208 692240 309240 692476
rect 308620 692156 309240 692240
rect 308620 691920 308652 692156
rect 308888 691920 308972 692156
rect 309208 691920 309240 692156
rect 344620 692240 344652 692476
rect 344888 692240 344972 692476
rect 345208 692240 345240 692476
rect 344620 692156 345240 692240
rect 344620 691920 344652 692156
rect 344888 691920 344972 692156
rect 345208 691920 345240 692156
rect 380620 692240 380652 692476
rect 380888 692240 380972 692476
rect 381208 692240 381240 692476
rect 380620 692156 381240 692240
rect 380620 691920 380652 692156
rect 380888 691920 380972 692156
rect 381208 691920 381240 692156
rect 416620 692240 416652 692476
rect 416888 692240 416972 692476
rect 417208 692240 417240 692476
rect 416620 692156 417240 692240
rect 416620 691920 416652 692156
rect 416888 691920 416972 692156
rect 417208 691920 417240 692156
rect 452620 692240 452652 692476
rect 452888 692240 452972 692476
rect 453208 692240 453240 692476
rect 452620 692156 453240 692240
rect 452620 691920 452652 692156
rect 452888 691920 452972 692156
rect 453208 691920 453240 692156
rect 488620 692240 488652 692476
rect 488888 692240 488972 692476
rect 489208 692240 489240 692476
rect 488620 692156 489240 692240
rect 488620 691920 488652 692156
rect 488888 691920 488972 692156
rect 489208 691920 489240 692156
rect 524620 692240 524652 692476
rect 524888 692240 524972 692476
rect 525208 692240 525240 692476
rect 524620 692156 525240 692240
rect 524620 691920 524652 692156
rect 524888 691920 524972 692156
rect 525208 691920 525240 692156
rect 560620 692240 560652 692476
rect 560888 692240 560972 692476
rect 561208 692240 561240 692476
rect 560620 692156 561240 692240
rect 560620 691920 560652 692156
rect 560888 691920 560972 692156
rect 561208 691920 561240 692156
rect 570260 692240 570292 692476
rect 570528 692240 570612 692476
rect 570848 692240 570880 692476
rect 570260 692156 570880 692240
rect 570260 691920 570292 692156
rect 570528 691920 570612 692156
rect 570848 691920 570880 692156
rect 7844 687138 7876 687374
rect 8112 687138 8196 687374
rect 8432 687138 8464 687374
rect 7844 687054 8464 687138
rect 7844 686818 7876 687054
rect 8112 686818 8196 687054
rect 8432 686818 8464 687054
rect 38000 687138 38032 687374
rect 38268 687138 38352 687374
rect 38588 687138 38620 687374
rect 38000 687054 38620 687138
rect 38000 686818 38032 687054
rect 38268 686818 38352 687054
rect 38588 686818 38620 687054
rect 74000 687138 74032 687374
rect 74268 687138 74352 687374
rect 74588 687138 74620 687374
rect 74000 687054 74620 687138
rect 74000 686818 74032 687054
rect 74268 686818 74352 687054
rect 74588 686818 74620 687054
rect 110000 687138 110032 687374
rect 110268 687138 110352 687374
rect 110588 687138 110620 687374
rect 110000 687054 110620 687138
rect 110000 686818 110032 687054
rect 110268 686818 110352 687054
rect 110588 686818 110620 687054
rect 146000 687138 146032 687374
rect 146268 687138 146352 687374
rect 146588 687138 146620 687374
rect 146000 687054 146620 687138
rect 146000 686818 146032 687054
rect 146268 686818 146352 687054
rect 146588 686818 146620 687054
rect 182000 687138 182032 687374
rect 182268 687138 182352 687374
rect 182588 687138 182620 687374
rect 182000 687054 182620 687138
rect 182000 686818 182032 687054
rect 182268 686818 182352 687054
rect 182588 686818 182620 687054
rect 218000 687138 218032 687374
rect 218268 687138 218352 687374
rect 218588 687138 218620 687374
rect 218000 687054 218620 687138
rect 218000 686818 218032 687054
rect 218268 686818 218352 687054
rect 218588 686818 218620 687054
rect 254000 687138 254032 687374
rect 254268 687138 254352 687374
rect 254588 687138 254620 687374
rect 254000 687054 254620 687138
rect 254000 686818 254032 687054
rect 254268 686818 254352 687054
rect 254588 686818 254620 687054
rect 290000 687138 290032 687374
rect 290268 687138 290352 687374
rect 290588 687138 290620 687374
rect 290000 687054 290620 687138
rect 290000 686818 290032 687054
rect 290268 686818 290352 687054
rect 290588 686818 290620 687054
rect 326000 687138 326032 687374
rect 326268 687138 326352 687374
rect 326588 687138 326620 687374
rect 326000 687054 326620 687138
rect 326000 686818 326032 687054
rect 326268 686818 326352 687054
rect 326588 686818 326620 687054
rect 362000 687138 362032 687374
rect 362268 687138 362352 687374
rect 362588 687138 362620 687374
rect 362000 687054 362620 687138
rect 362000 686818 362032 687054
rect 362268 686818 362352 687054
rect 362588 686818 362620 687054
rect 398000 687138 398032 687374
rect 398268 687138 398352 687374
rect 398588 687138 398620 687374
rect 398000 687054 398620 687138
rect 398000 686818 398032 687054
rect 398268 686818 398352 687054
rect 398588 686818 398620 687054
rect 434000 687138 434032 687374
rect 434268 687138 434352 687374
rect 434588 687138 434620 687374
rect 434000 687054 434620 687138
rect 434000 686818 434032 687054
rect 434268 686818 434352 687054
rect 434588 686818 434620 687054
rect 470000 687138 470032 687374
rect 470268 687138 470352 687374
rect 470588 687138 470620 687374
rect 470000 687054 470620 687138
rect 470000 686818 470032 687054
rect 470268 686818 470352 687054
rect 470588 686818 470620 687054
rect 506000 687138 506032 687374
rect 506268 687138 506352 687374
rect 506588 687138 506620 687374
rect 506000 687054 506620 687138
rect 506000 686818 506032 687054
rect 506268 686818 506352 687054
rect 506588 686818 506620 687054
rect 542000 687138 542032 687374
rect 542268 687138 542352 687374
rect 542588 687138 542620 687374
rect 542000 687054 542620 687138
rect 542000 686818 542032 687054
rect 542268 686818 542352 687054
rect 542588 686818 542620 687054
rect 571500 687138 571532 687374
rect 571768 687138 571852 687374
rect 572088 687138 572120 687374
rect 571500 687054 572120 687138
rect 571500 686818 571532 687054
rect 571768 686818 571852 687054
rect 572088 686818 572120 687054
rect -2006 683418 -1974 683654
rect -1738 683418 -1654 683654
rect -1418 683418 -1386 683654
rect -2006 683334 -1386 683418
rect -2006 683098 -1974 683334
rect -1738 683098 -1654 683334
rect -1418 683098 -1386 683334
rect 9084 683418 9116 683654
rect 9352 683418 9436 683654
rect 9672 683418 9704 683654
rect 9084 683334 9704 683418
rect 9084 683098 9116 683334
rect 9352 683098 9436 683334
rect 9672 683098 9704 683334
rect 56620 683418 56652 683654
rect 56888 683418 56972 683654
rect 57208 683418 57240 683654
rect 56620 683334 57240 683418
rect 56620 683098 56652 683334
rect 56888 683098 56972 683334
rect 57208 683098 57240 683334
rect 92620 683418 92652 683654
rect 92888 683418 92972 683654
rect 93208 683418 93240 683654
rect 92620 683334 93240 683418
rect 92620 683098 92652 683334
rect 92888 683098 92972 683334
rect 93208 683098 93240 683334
rect 128620 683418 128652 683654
rect 128888 683418 128972 683654
rect 129208 683418 129240 683654
rect 128620 683334 129240 683418
rect 128620 683098 128652 683334
rect 128888 683098 128972 683334
rect 129208 683098 129240 683334
rect 164620 683418 164652 683654
rect 164888 683418 164972 683654
rect 165208 683418 165240 683654
rect 164620 683334 165240 683418
rect 164620 683098 164652 683334
rect 164888 683098 164972 683334
rect 165208 683098 165240 683334
rect 200620 683418 200652 683654
rect 200888 683418 200972 683654
rect 201208 683418 201240 683654
rect 200620 683334 201240 683418
rect 200620 683098 200652 683334
rect 200888 683098 200972 683334
rect 201208 683098 201240 683334
rect 236620 683418 236652 683654
rect 236888 683418 236972 683654
rect 237208 683418 237240 683654
rect 236620 683334 237240 683418
rect 236620 683098 236652 683334
rect 236888 683098 236972 683334
rect 237208 683098 237240 683334
rect 272620 683418 272652 683654
rect 272888 683418 272972 683654
rect 273208 683418 273240 683654
rect 272620 683334 273240 683418
rect 272620 683098 272652 683334
rect 272888 683098 272972 683334
rect 273208 683098 273240 683334
rect 308620 683418 308652 683654
rect 308888 683418 308972 683654
rect 309208 683418 309240 683654
rect 308620 683334 309240 683418
rect 308620 683098 308652 683334
rect 308888 683098 308972 683334
rect 309208 683098 309240 683334
rect 344620 683418 344652 683654
rect 344888 683418 344972 683654
rect 345208 683418 345240 683654
rect 344620 683334 345240 683418
rect 344620 683098 344652 683334
rect 344888 683098 344972 683334
rect 345208 683098 345240 683334
rect 380620 683418 380652 683654
rect 380888 683418 380972 683654
rect 381208 683418 381240 683654
rect 380620 683334 381240 683418
rect 380620 683098 380652 683334
rect 380888 683098 380972 683334
rect 381208 683098 381240 683334
rect 416620 683418 416652 683654
rect 416888 683418 416972 683654
rect 417208 683418 417240 683654
rect 416620 683334 417240 683418
rect 416620 683098 416652 683334
rect 416888 683098 416972 683334
rect 417208 683098 417240 683334
rect 452620 683418 452652 683654
rect 452888 683418 452972 683654
rect 453208 683418 453240 683654
rect 452620 683334 453240 683418
rect 452620 683098 452652 683334
rect 452888 683098 452972 683334
rect 453208 683098 453240 683334
rect 488620 683418 488652 683654
rect 488888 683418 488972 683654
rect 489208 683418 489240 683654
rect 488620 683334 489240 683418
rect 488620 683098 488652 683334
rect 488888 683098 488972 683334
rect 489208 683098 489240 683334
rect 524620 683418 524652 683654
rect 524888 683418 524972 683654
rect 525208 683418 525240 683654
rect 524620 683334 525240 683418
rect 524620 683098 524652 683334
rect 524888 683098 524972 683334
rect 525208 683098 525240 683334
rect 560620 683418 560652 683654
rect 560888 683418 560972 683654
rect 561208 683418 561240 683654
rect 560620 683334 561240 683418
rect 560620 683098 560652 683334
rect 560888 683098 560972 683334
rect 561208 683098 561240 683334
rect 570260 683418 570292 683654
rect 570528 683418 570612 683654
rect 570848 683418 570880 683654
rect 570260 683334 570880 683418
rect 570260 683098 570292 683334
rect 570528 683098 570612 683334
rect 570848 683098 570880 683334
rect -2006 643654 -1386 683098
rect 580594 662254 581214 719832
rect 600860 720388 601480 720420
rect 600860 720152 600892 720388
rect 601128 720152 601212 720388
rect 601448 720152 601480 720388
rect 600860 720068 601480 720152
rect 600860 719832 600892 720068
rect 601128 719832 601212 720068
rect 601448 719832 601480 720068
rect 597750 717278 598370 717310
rect 597750 717042 597782 717278
rect 598018 717042 598102 717278
rect 598338 717042 598370 717278
rect 597750 716958 598370 717042
rect 597750 716722 597782 716958
rect 598018 716722 598102 716958
rect 598338 716722 598370 716958
rect 594640 714168 595260 714200
rect 594640 713932 594672 714168
rect 594908 713932 594992 714168
rect 595228 713932 595260 714168
rect 594640 713848 595260 713932
rect 594640 713612 594672 713848
rect 594908 713612 594992 713848
rect 595228 713612 595260 713848
rect 591530 711058 592150 711090
rect 591530 710822 591562 711058
rect 591798 710822 591882 711058
rect 592118 710822 592150 711058
rect 591530 710738 592150 710822
rect 591530 710502 591562 710738
rect 591798 710502 591882 710738
rect 592118 710502 592150 710738
rect 588420 707948 589040 707980
rect 588420 707712 588452 707948
rect 588688 707712 588772 707948
rect 589008 707712 589040 707948
rect 588420 707628 589040 707712
rect 588420 707392 588452 707628
rect 588688 707392 588772 707628
rect 589008 707392 589040 707628
rect 580594 662018 580626 662254
rect 580862 662018 580946 662254
rect 581182 662018 581214 662254
rect 580594 661934 581214 662018
rect 580594 661698 580626 661934
rect 580862 661698 580946 661934
rect 581182 661698 581214 661934
rect 7844 647138 7876 647374
rect 8112 647138 8196 647374
rect 8432 647138 8464 647374
rect 7844 647054 8464 647138
rect 7844 646818 7876 647054
rect 8112 646818 8196 647054
rect 8432 646818 8464 647054
rect 38000 647138 38032 647374
rect 38268 647138 38352 647374
rect 38588 647138 38620 647374
rect 38000 647054 38620 647138
rect 38000 646818 38032 647054
rect 38268 646818 38352 647054
rect 38588 646818 38620 647054
rect 74000 647138 74032 647374
rect 74268 647138 74352 647374
rect 74588 647138 74620 647374
rect 74000 647054 74620 647138
rect 74000 646818 74032 647054
rect 74268 646818 74352 647054
rect 74588 646818 74620 647054
rect 110000 647138 110032 647374
rect 110268 647138 110352 647374
rect 110588 647138 110620 647374
rect 110000 647054 110620 647138
rect 110000 646818 110032 647054
rect 110268 646818 110352 647054
rect 110588 646818 110620 647054
rect 146000 647138 146032 647374
rect 146268 647138 146352 647374
rect 146588 647138 146620 647374
rect 146000 647054 146620 647138
rect 146000 646818 146032 647054
rect 146268 646818 146352 647054
rect 146588 646818 146620 647054
rect 182000 647138 182032 647374
rect 182268 647138 182352 647374
rect 182588 647138 182620 647374
rect 182000 647054 182620 647138
rect 182000 646818 182032 647054
rect 182268 646818 182352 647054
rect 182588 646818 182620 647054
rect 218000 647138 218032 647374
rect 218268 647138 218352 647374
rect 218588 647138 218620 647374
rect 218000 647054 218620 647138
rect 218000 646818 218032 647054
rect 218268 646818 218352 647054
rect 218588 646818 218620 647054
rect 254000 647138 254032 647374
rect 254268 647138 254352 647374
rect 254588 647138 254620 647374
rect 254000 647054 254620 647138
rect 254000 646818 254032 647054
rect 254268 646818 254352 647054
rect 254588 646818 254620 647054
rect 290000 647138 290032 647374
rect 290268 647138 290352 647374
rect 290588 647138 290620 647374
rect 290000 647054 290620 647138
rect 290000 646818 290032 647054
rect 290268 646818 290352 647054
rect 290588 646818 290620 647054
rect 326000 647138 326032 647374
rect 326268 647138 326352 647374
rect 326588 647138 326620 647374
rect 326000 647054 326620 647138
rect 326000 646818 326032 647054
rect 326268 646818 326352 647054
rect 326588 646818 326620 647054
rect 362000 647138 362032 647374
rect 362268 647138 362352 647374
rect 362588 647138 362620 647374
rect 362000 647054 362620 647138
rect 362000 646818 362032 647054
rect 362268 646818 362352 647054
rect 362588 646818 362620 647054
rect 398000 647138 398032 647374
rect 398268 647138 398352 647374
rect 398588 647138 398620 647374
rect 398000 647054 398620 647138
rect 398000 646818 398032 647054
rect 398268 646818 398352 647054
rect 398588 646818 398620 647054
rect 434000 647138 434032 647374
rect 434268 647138 434352 647374
rect 434588 647138 434620 647374
rect 434000 647054 434620 647138
rect 434000 646818 434032 647054
rect 434268 646818 434352 647054
rect 434588 646818 434620 647054
rect 470000 647138 470032 647374
rect 470268 647138 470352 647374
rect 470588 647138 470620 647374
rect 470000 647054 470620 647138
rect 470000 646818 470032 647054
rect 470268 646818 470352 647054
rect 470588 646818 470620 647054
rect 506000 647138 506032 647374
rect 506268 647138 506352 647374
rect 506588 647138 506620 647374
rect 506000 647054 506620 647138
rect 506000 646818 506032 647054
rect 506268 646818 506352 647054
rect 506588 646818 506620 647054
rect 542000 647138 542032 647374
rect 542268 647138 542352 647374
rect 542588 647138 542620 647374
rect 542000 647054 542620 647138
rect 542000 646818 542032 647054
rect 542268 646818 542352 647054
rect 542588 646818 542620 647054
rect 571500 647138 571532 647374
rect 571768 647138 571852 647374
rect 572088 647138 572120 647374
rect 571500 647054 572120 647138
rect 571500 646818 571532 647054
rect 571768 646818 571852 647054
rect 572088 646818 572120 647054
rect -2006 643418 -1974 643654
rect -1738 643418 -1654 643654
rect -1418 643418 -1386 643654
rect -2006 643334 -1386 643418
rect -2006 643098 -1974 643334
rect -1738 643098 -1654 643334
rect -1418 643098 -1386 643334
rect 9084 643418 9116 643654
rect 9352 643418 9436 643654
rect 9672 643418 9704 643654
rect 9084 643334 9704 643418
rect 9084 643098 9116 643334
rect 9352 643098 9436 643334
rect 9672 643098 9704 643334
rect 56620 643418 56652 643654
rect 56888 643418 56972 643654
rect 57208 643418 57240 643654
rect 56620 643334 57240 643418
rect 56620 643098 56652 643334
rect 56888 643098 56972 643334
rect 57208 643098 57240 643334
rect 92620 643418 92652 643654
rect 92888 643418 92972 643654
rect 93208 643418 93240 643654
rect 92620 643334 93240 643418
rect 92620 643098 92652 643334
rect 92888 643098 92972 643334
rect 93208 643098 93240 643334
rect 128620 643418 128652 643654
rect 128888 643418 128972 643654
rect 129208 643418 129240 643654
rect 128620 643334 129240 643418
rect 128620 643098 128652 643334
rect 128888 643098 128972 643334
rect 129208 643098 129240 643334
rect 164620 643418 164652 643654
rect 164888 643418 164972 643654
rect 165208 643418 165240 643654
rect 164620 643334 165240 643418
rect 164620 643098 164652 643334
rect 164888 643098 164972 643334
rect 165208 643098 165240 643334
rect 200620 643418 200652 643654
rect 200888 643418 200972 643654
rect 201208 643418 201240 643654
rect 200620 643334 201240 643418
rect 200620 643098 200652 643334
rect 200888 643098 200972 643334
rect 201208 643098 201240 643334
rect 236620 643418 236652 643654
rect 236888 643418 236972 643654
rect 237208 643418 237240 643654
rect 236620 643334 237240 643418
rect 236620 643098 236652 643334
rect 236888 643098 236972 643334
rect 237208 643098 237240 643334
rect 272620 643418 272652 643654
rect 272888 643418 272972 643654
rect 273208 643418 273240 643654
rect 272620 643334 273240 643418
rect 272620 643098 272652 643334
rect 272888 643098 272972 643334
rect 273208 643098 273240 643334
rect 308620 643418 308652 643654
rect 308888 643418 308972 643654
rect 309208 643418 309240 643654
rect 308620 643334 309240 643418
rect 308620 643098 308652 643334
rect 308888 643098 308972 643334
rect 309208 643098 309240 643334
rect 344620 643418 344652 643654
rect 344888 643418 344972 643654
rect 345208 643418 345240 643654
rect 344620 643334 345240 643418
rect 344620 643098 344652 643334
rect 344888 643098 344972 643334
rect 345208 643098 345240 643334
rect 380620 643418 380652 643654
rect 380888 643418 380972 643654
rect 381208 643418 381240 643654
rect 380620 643334 381240 643418
rect 380620 643098 380652 643334
rect 380888 643098 380972 643334
rect 381208 643098 381240 643334
rect 416620 643418 416652 643654
rect 416888 643418 416972 643654
rect 417208 643418 417240 643654
rect 416620 643334 417240 643418
rect 416620 643098 416652 643334
rect 416888 643098 416972 643334
rect 417208 643098 417240 643334
rect 452620 643418 452652 643654
rect 452888 643418 452972 643654
rect 453208 643418 453240 643654
rect 452620 643334 453240 643418
rect 452620 643098 452652 643334
rect 452888 643098 452972 643334
rect 453208 643098 453240 643334
rect 488620 643418 488652 643654
rect 488888 643418 488972 643654
rect 489208 643418 489240 643654
rect 488620 643334 489240 643418
rect 488620 643098 488652 643334
rect 488888 643098 488972 643334
rect 489208 643098 489240 643334
rect 524620 643418 524652 643654
rect 524888 643418 524972 643654
rect 525208 643418 525240 643654
rect 524620 643334 525240 643418
rect 524620 643098 524652 643334
rect 524888 643098 524972 643334
rect 525208 643098 525240 643334
rect 560620 643418 560652 643654
rect 560888 643418 560972 643654
rect 561208 643418 561240 643654
rect 560620 643334 561240 643418
rect 560620 643098 560652 643334
rect 560888 643098 560972 643334
rect 561208 643098 561240 643334
rect 570260 643418 570292 643654
rect 570528 643418 570612 643654
rect 570848 643418 570880 643654
rect 570260 643334 570880 643418
rect 570260 643098 570292 643334
rect 570528 643098 570612 643334
rect 570848 643098 570880 643334
rect -2006 603654 -1386 643098
rect 580594 622254 581214 661698
rect 580594 622018 580626 622254
rect 580862 622018 580946 622254
rect 581182 622018 581214 622254
rect 580594 621934 581214 622018
rect 580594 621698 580626 621934
rect 580862 621698 580946 621934
rect 581182 621698 581214 621934
rect 7844 607138 7876 607374
rect 8112 607138 8196 607374
rect 8432 607138 8464 607374
rect 7844 607054 8464 607138
rect 7844 606818 7876 607054
rect 8112 606818 8196 607054
rect 8432 606818 8464 607054
rect 38000 607138 38032 607374
rect 38268 607138 38352 607374
rect 38588 607138 38620 607374
rect 38000 607054 38620 607138
rect 38000 606818 38032 607054
rect 38268 606818 38352 607054
rect 38588 606818 38620 607054
rect 74000 607138 74032 607374
rect 74268 607138 74352 607374
rect 74588 607138 74620 607374
rect 74000 607054 74620 607138
rect 74000 606818 74032 607054
rect 74268 606818 74352 607054
rect 74588 606818 74620 607054
rect 110000 607138 110032 607374
rect 110268 607138 110352 607374
rect 110588 607138 110620 607374
rect 110000 607054 110620 607138
rect 110000 606818 110032 607054
rect 110268 606818 110352 607054
rect 110588 606818 110620 607054
rect 146000 607138 146032 607374
rect 146268 607138 146352 607374
rect 146588 607138 146620 607374
rect 146000 607054 146620 607138
rect 146000 606818 146032 607054
rect 146268 606818 146352 607054
rect 146588 606818 146620 607054
rect 182000 607138 182032 607374
rect 182268 607138 182352 607374
rect 182588 607138 182620 607374
rect 182000 607054 182620 607138
rect 182000 606818 182032 607054
rect 182268 606818 182352 607054
rect 182588 606818 182620 607054
rect 218000 607138 218032 607374
rect 218268 607138 218352 607374
rect 218588 607138 218620 607374
rect 218000 607054 218620 607138
rect 218000 606818 218032 607054
rect 218268 606818 218352 607054
rect 218588 606818 218620 607054
rect 254000 607138 254032 607374
rect 254268 607138 254352 607374
rect 254588 607138 254620 607374
rect 254000 607054 254620 607138
rect 254000 606818 254032 607054
rect 254268 606818 254352 607054
rect 254588 606818 254620 607054
rect 290000 607138 290032 607374
rect 290268 607138 290352 607374
rect 290588 607138 290620 607374
rect 290000 607054 290620 607138
rect 290000 606818 290032 607054
rect 290268 606818 290352 607054
rect 290588 606818 290620 607054
rect 326000 607138 326032 607374
rect 326268 607138 326352 607374
rect 326588 607138 326620 607374
rect 326000 607054 326620 607138
rect 326000 606818 326032 607054
rect 326268 606818 326352 607054
rect 326588 606818 326620 607054
rect 362000 607138 362032 607374
rect 362268 607138 362352 607374
rect 362588 607138 362620 607374
rect 362000 607054 362620 607138
rect 362000 606818 362032 607054
rect 362268 606818 362352 607054
rect 362588 606818 362620 607054
rect 398000 607138 398032 607374
rect 398268 607138 398352 607374
rect 398588 607138 398620 607374
rect 398000 607054 398620 607138
rect 398000 606818 398032 607054
rect 398268 606818 398352 607054
rect 398588 606818 398620 607054
rect 434000 607138 434032 607374
rect 434268 607138 434352 607374
rect 434588 607138 434620 607374
rect 434000 607054 434620 607138
rect 434000 606818 434032 607054
rect 434268 606818 434352 607054
rect 434588 606818 434620 607054
rect 470000 607138 470032 607374
rect 470268 607138 470352 607374
rect 470588 607138 470620 607374
rect 470000 607054 470620 607138
rect 470000 606818 470032 607054
rect 470268 606818 470352 607054
rect 470588 606818 470620 607054
rect 506000 607138 506032 607374
rect 506268 607138 506352 607374
rect 506588 607138 506620 607374
rect 506000 607054 506620 607138
rect 506000 606818 506032 607054
rect 506268 606818 506352 607054
rect 506588 606818 506620 607054
rect 542000 607138 542032 607374
rect 542268 607138 542352 607374
rect 542588 607138 542620 607374
rect 542000 607054 542620 607138
rect 542000 606818 542032 607054
rect 542268 606818 542352 607054
rect 542588 606818 542620 607054
rect 571500 607138 571532 607374
rect 571768 607138 571852 607374
rect 572088 607138 572120 607374
rect 571500 607054 572120 607138
rect 571500 606818 571532 607054
rect 571768 606818 571852 607054
rect 572088 606818 572120 607054
rect -2006 603418 -1974 603654
rect -1738 603418 -1654 603654
rect -1418 603418 -1386 603654
rect -2006 603334 -1386 603418
rect -2006 603098 -1974 603334
rect -1738 603098 -1654 603334
rect -1418 603098 -1386 603334
rect 9084 603418 9116 603654
rect 9352 603418 9436 603654
rect 9672 603418 9704 603654
rect 9084 603334 9704 603418
rect 9084 603098 9116 603334
rect 9352 603098 9436 603334
rect 9672 603098 9704 603334
rect 56620 603418 56652 603654
rect 56888 603418 56972 603654
rect 57208 603418 57240 603654
rect 56620 603334 57240 603418
rect 56620 603098 56652 603334
rect 56888 603098 56972 603334
rect 57208 603098 57240 603334
rect 92620 603418 92652 603654
rect 92888 603418 92972 603654
rect 93208 603418 93240 603654
rect 92620 603334 93240 603418
rect 92620 603098 92652 603334
rect 92888 603098 92972 603334
rect 93208 603098 93240 603334
rect 128620 603418 128652 603654
rect 128888 603418 128972 603654
rect 129208 603418 129240 603654
rect 128620 603334 129240 603418
rect 128620 603098 128652 603334
rect 128888 603098 128972 603334
rect 129208 603098 129240 603334
rect 164620 603418 164652 603654
rect 164888 603418 164972 603654
rect 165208 603418 165240 603654
rect 164620 603334 165240 603418
rect 164620 603098 164652 603334
rect 164888 603098 164972 603334
rect 165208 603098 165240 603334
rect 200620 603418 200652 603654
rect 200888 603418 200972 603654
rect 201208 603418 201240 603654
rect 200620 603334 201240 603418
rect 200620 603098 200652 603334
rect 200888 603098 200972 603334
rect 201208 603098 201240 603334
rect 236620 603418 236652 603654
rect 236888 603418 236972 603654
rect 237208 603418 237240 603654
rect 236620 603334 237240 603418
rect 236620 603098 236652 603334
rect 236888 603098 236972 603334
rect 237208 603098 237240 603334
rect 272620 603418 272652 603654
rect 272888 603418 272972 603654
rect 273208 603418 273240 603654
rect 272620 603334 273240 603418
rect 272620 603098 272652 603334
rect 272888 603098 272972 603334
rect 273208 603098 273240 603334
rect 308620 603418 308652 603654
rect 308888 603418 308972 603654
rect 309208 603418 309240 603654
rect 308620 603334 309240 603418
rect 308620 603098 308652 603334
rect 308888 603098 308972 603334
rect 309208 603098 309240 603334
rect 344620 603418 344652 603654
rect 344888 603418 344972 603654
rect 345208 603418 345240 603654
rect 344620 603334 345240 603418
rect 344620 603098 344652 603334
rect 344888 603098 344972 603334
rect 345208 603098 345240 603334
rect 380620 603418 380652 603654
rect 380888 603418 380972 603654
rect 381208 603418 381240 603654
rect 380620 603334 381240 603418
rect 380620 603098 380652 603334
rect 380888 603098 380972 603334
rect 381208 603098 381240 603334
rect 416620 603418 416652 603654
rect 416888 603418 416972 603654
rect 417208 603418 417240 603654
rect 416620 603334 417240 603418
rect 416620 603098 416652 603334
rect 416888 603098 416972 603334
rect 417208 603098 417240 603334
rect 452620 603418 452652 603654
rect 452888 603418 452972 603654
rect 453208 603418 453240 603654
rect 452620 603334 453240 603418
rect 452620 603098 452652 603334
rect 452888 603098 452972 603334
rect 453208 603098 453240 603334
rect 488620 603418 488652 603654
rect 488888 603418 488972 603654
rect 489208 603418 489240 603654
rect 488620 603334 489240 603418
rect 488620 603098 488652 603334
rect 488888 603098 488972 603334
rect 489208 603098 489240 603334
rect 524620 603418 524652 603654
rect 524888 603418 524972 603654
rect 525208 603418 525240 603654
rect 524620 603334 525240 603418
rect 524620 603098 524652 603334
rect 524888 603098 524972 603334
rect 525208 603098 525240 603334
rect 560620 603418 560652 603654
rect 560888 603418 560972 603654
rect 561208 603418 561240 603654
rect 560620 603334 561240 603418
rect 560620 603098 560652 603334
rect 560888 603098 560972 603334
rect 561208 603098 561240 603334
rect 570260 603418 570292 603654
rect 570528 603418 570612 603654
rect 570848 603418 570880 603654
rect 570260 603334 570880 603418
rect 570260 603098 570292 603334
rect 570528 603098 570612 603334
rect 570848 603098 570880 603334
rect -2006 563654 -1386 603098
rect 580594 582254 581214 621698
rect 580594 582018 580626 582254
rect 580862 582018 580946 582254
rect 581182 582018 581214 582254
rect 580594 581934 581214 582018
rect 580594 581698 580626 581934
rect 580862 581698 580946 581934
rect 581182 581698 581214 581934
rect 7844 567138 7876 567374
rect 8112 567138 8196 567374
rect 8432 567138 8464 567374
rect 7844 567054 8464 567138
rect 7844 566818 7876 567054
rect 8112 566818 8196 567054
rect 8432 566818 8464 567054
rect 38000 567138 38032 567374
rect 38268 567138 38352 567374
rect 38588 567138 38620 567374
rect 38000 567054 38620 567138
rect 38000 566818 38032 567054
rect 38268 566818 38352 567054
rect 38588 566818 38620 567054
rect 74000 567138 74032 567374
rect 74268 567138 74352 567374
rect 74588 567138 74620 567374
rect 74000 567054 74620 567138
rect 74000 566818 74032 567054
rect 74268 566818 74352 567054
rect 74588 566818 74620 567054
rect 110000 567138 110032 567374
rect 110268 567138 110352 567374
rect 110588 567138 110620 567374
rect 110000 567054 110620 567138
rect 110000 566818 110032 567054
rect 110268 566818 110352 567054
rect 110588 566818 110620 567054
rect 146000 567138 146032 567374
rect 146268 567138 146352 567374
rect 146588 567138 146620 567374
rect 146000 567054 146620 567138
rect 146000 566818 146032 567054
rect 146268 566818 146352 567054
rect 146588 566818 146620 567054
rect 182000 567138 182032 567374
rect 182268 567138 182352 567374
rect 182588 567138 182620 567374
rect 182000 567054 182620 567138
rect 182000 566818 182032 567054
rect 182268 566818 182352 567054
rect 182588 566818 182620 567054
rect 218000 567138 218032 567374
rect 218268 567138 218352 567374
rect 218588 567138 218620 567374
rect 218000 567054 218620 567138
rect 218000 566818 218032 567054
rect 218268 566818 218352 567054
rect 218588 566818 218620 567054
rect 254000 567138 254032 567374
rect 254268 567138 254352 567374
rect 254588 567138 254620 567374
rect 254000 567054 254620 567138
rect 254000 566818 254032 567054
rect 254268 566818 254352 567054
rect 254588 566818 254620 567054
rect 290000 567138 290032 567374
rect 290268 567138 290352 567374
rect 290588 567138 290620 567374
rect 290000 567054 290620 567138
rect 290000 566818 290032 567054
rect 290268 566818 290352 567054
rect 290588 566818 290620 567054
rect 326000 567138 326032 567374
rect 326268 567138 326352 567374
rect 326588 567138 326620 567374
rect 326000 567054 326620 567138
rect 326000 566818 326032 567054
rect 326268 566818 326352 567054
rect 326588 566818 326620 567054
rect 362000 567138 362032 567374
rect 362268 567138 362352 567374
rect 362588 567138 362620 567374
rect 362000 567054 362620 567138
rect 362000 566818 362032 567054
rect 362268 566818 362352 567054
rect 362588 566818 362620 567054
rect 398000 567138 398032 567374
rect 398268 567138 398352 567374
rect 398588 567138 398620 567374
rect 398000 567054 398620 567138
rect 398000 566818 398032 567054
rect 398268 566818 398352 567054
rect 398588 566818 398620 567054
rect 434000 567138 434032 567374
rect 434268 567138 434352 567374
rect 434588 567138 434620 567374
rect 434000 567054 434620 567138
rect 434000 566818 434032 567054
rect 434268 566818 434352 567054
rect 434588 566818 434620 567054
rect 470000 567138 470032 567374
rect 470268 567138 470352 567374
rect 470588 567138 470620 567374
rect 470000 567054 470620 567138
rect 470000 566818 470032 567054
rect 470268 566818 470352 567054
rect 470588 566818 470620 567054
rect 506000 567138 506032 567374
rect 506268 567138 506352 567374
rect 506588 567138 506620 567374
rect 506000 567054 506620 567138
rect 506000 566818 506032 567054
rect 506268 566818 506352 567054
rect 506588 566818 506620 567054
rect 542000 567138 542032 567374
rect 542268 567138 542352 567374
rect 542588 567138 542620 567374
rect 542000 567054 542620 567138
rect 542000 566818 542032 567054
rect 542268 566818 542352 567054
rect 542588 566818 542620 567054
rect 571500 567138 571532 567374
rect 571768 567138 571852 567374
rect 572088 567138 572120 567374
rect 571500 567054 572120 567138
rect 571500 566818 571532 567054
rect 571768 566818 571852 567054
rect 572088 566818 572120 567054
rect -2006 563418 -1974 563654
rect -1738 563418 -1654 563654
rect -1418 563418 -1386 563654
rect -2006 563334 -1386 563418
rect -2006 563098 -1974 563334
rect -1738 563098 -1654 563334
rect -1418 563098 -1386 563334
rect 9084 563418 9116 563654
rect 9352 563418 9436 563654
rect 9672 563418 9704 563654
rect 9084 563334 9704 563418
rect 9084 563098 9116 563334
rect 9352 563098 9436 563334
rect 9672 563098 9704 563334
rect 56620 563418 56652 563654
rect 56888 563418 56972 563654
rect 57208 563418 57240 563654
rect 56620 563334 57240 563418
rect 56620 563098 56652 563334
rect 56888 563098 56972 563334
rect 57208 563098 57240 563334
rect 92620 563418 92652 563654
rect 92888 563418 92972 563654
rect 93208 563418 93240 563654
rect 92620 563334 93240 563418
rect 92620 563098 92652 563334
rect 92888 563098 92972 563334
rect 93208 563098 93240 563334
rect 128620 563418 128652 563654
rect 128888 563418 128972 563654
rect 129208 563418 129240 563654
rect 128620 563334 129240 563418
rect 128620 563098 128652 563334
rect 128888 563098 128972 563334
rect 129208 563098 129240 563334
rect 164620 563418 164652 563654
rect 164888 563418 164972 563654
rect 165208 563418 165240 563654
rect 164620 563334 165240 563418
rect 164620 563098 164652 563334
rect 164888 563098 164972 563334
rect 165208 563098 165240 563334
rect 200620 563418 200652 563654
rect 200888 563418 200972 563654
rect 201208 563418 201240 563654
rect 200620 563334 201240 563418
rect 200620 563098 200652 563334
rect 200888 563098 200972 563334
rect 201208 563098 201240 563334
rect 236620 563418 236652 563654
rect 236888 563418 236972 563654
rect 237208 563418 237240 563654
rect 236620 563334 237240 563418
rect 236620 563098 236652 563334
rect 236888 563098 236972 563334
rect 237208 563098 237240 563334
rect 272620 563418 272652 563654
rect 272888 563418 272972 563654
rect 273208 563418 273240 563654
rect 272620 563334 273240 563418
rect 272620 563098 272652 563334
rect 272888 563098 272972 563334
rect 273208 563098 273240 563334
rect 308620 563418 308652 563654
rect 308888 563418 308972 563654
rect 309208 563418 309240 563654
rect 308620 563334 309240 563418
rect 308620 563098 308652 563334
rect 308888 563098 308972 563334
rect 309208 563098 309240 563334
rect 344620 563418 344652 563654
rect 344888 563418 344972 563654
rect 345208 563418 345240 563654
rect 344620 563334 345240 563418
rect 344620 563098 344652 563334
rect 344888 563098 344972 563334
rect 345208 563098 345240 563334
rect 380620 563418 380652 563654
rect 380888 563418 380972 563654
rect 381208 563418 381240 563654
rect 380620 563334 381240 563418
rect 380620 563098 380652 563334
rect 380888 563098 380972 563334
rect 381208 563098 381240 563334
rect 416620 563418 416652 563654
rect 416888 563418 416972 563654
rect 417208 563418 417240 563654
rect 416620 563334 417240 563418
rect 416620 563098 416652 563334
rect 416888 563098 416972 563334
rect 417208 563098 417240 563334
rect 452620 563418 452652 563654
rect 452888 563418 452972 563654
rect 453208 563418 453240 563654
rect 452620 563334 453240 563418
rect 452620 563098 452652 563334
rect 452888 563098 452972 563334
rect 453208 563098 453240 563334
rect 488620 563418 488652 563654
rect 488888 563418 488972 563654
rect 489208 563418 489240 563654
rect 488620 563334 489240 563418
rect 488620 563098 488652 563334
rect 488888 563098 488972 563334
rect 489208 563098 489240 563334
rect 524620 563418 524652 563654
rect 524888 563418 524972 563654
rect 525208 563418 525240 563654
rect 524620 563334 525240 563418
rect 524620 563098 524652 563334
rect 524888 563098 524972 563334
rect 525208 563098 525240 563334
rect 560620 563418 560652 563654
rect 560888 563418 560972 563654
rect 561208 563418 561240 563654
rect 560620 563334 561240 563418
rect 560620 563098 560652 563334
rect 560888 563098 560972 563334
rect 561208 563098 561240 563334
rect 570260 563418 570292 563654
rect 570528 563418 570612 563654
rect 570848 563418 570880 563654
rect 570260 563334 570880 563418
rect 570260 563098 570292 563334
rect 570528 563098 570612 563334
rect 570848 563098 570880 563334
rect -2006 523654 -1386 563098
rect 580594 542254 581214 581698
rect 580594 542018 580626 542254
rect 580862 542018 580946 542254
rect 581182 542018 581214 542254
rect 580594 541934 581214 542018
rect 580594 541698 580626 541934
rect 580862 541698 580946 541934
rect 581182 541698 581214 541934
rect 7844 527138 7876 527374
rect 8112 527138 8196 527374
rect 8432 527138 8464 527374
rect 7844 527054 8464 527138
rect 7844 526818 7876 527054
rect 8112 526818 8196 527054
rect 8432 526818 8464 527054
rect 38000 527138 38032 527374
rect 38268 527138 38352 527374
rect 38588 527138 38620 527374
rect 38000 527054 38620 527138
rect 38000 526818 38032 527054
rect 38268 526818 38352 527054
rect 38588 526818 38620 527054
rect 74000 527138 74032 527374
rect 74268 527138 74352 527374
rect 74588 527138 74620 527374
rect 74000 527054 74620 527138
rect 74000 526818 74032 527054
rect 74268 526818 74352 527054
rect 74588 526818 74620 527054
rect 110000 527138 110032 527374
rect 110268 527138 110352 527374
rect 110588 527138 110620 527374
rect 110000 527054 110620 527138
rect 110000 526818 110032 527054
rect 110268 526818 110352 527054
rect 110588 526818 110620 527054
rect 146000 527138 146032 527374
rect 146268 527138 146352 527374
rect 146588 527138 146620 527374
rect 146000 527054 146620 527138
rect 146000 526818 146032 527054
rect 146268 526818 146352 527054
rect 146588 526818 146620 527054
rect 182000 527138 182032 527374
rect 182268 527138 182352 527374
rect 182588 527138 182620 527374
rect 182000 527054 182620 527138
rect 182000 526818 182032 527054
rect 182268 526818 182352 527054
rect 182588 526818 182620 527054
rect 218000 527138 218032 527374
rect 218268 527138 218352 527374
rect 218588 527138 218620 527374
rect 218000 527054 218620 527138
rect 218000 526818 218032 527054
rect 218268 526818 218352 527054
rect 218588 526818 218620 527054
rect 254000 527138 254032 527374
rect 254268 527138 254352 527374
rect 254588 527138 254620 527374
rect 254000 527054 254620 527138
rect 254000 526818 254032 527054
rect 254268 526818 254352 527054
rect 254588 526818 254620 527054
rect 290000 527138 290032 527374
rect 290268 527138 290352 527374
rect 290588 527138 290620 527374
rect 290000 527054 290620 527138
rect 290000 526818 290032 527054
rect 290268 526818 290352 527054
rect 290588 526818 290620 527054
rect 326000 527138 326032 527374
rect 326268 527138 326352 527374
rect 326588 527138 326620 527374
rect 326000 527054 326620 527138
rect 326000 526818 326032 527054
rect 326268 526818 326352 527054
rect 326588 526818 326620 527054
rect 362000 527138 362032 527374
rect 362268 527138 362352 527374
rect 362588 527138 362620 527374
rect 362000 527054 362620 527138
rect 362000 526818 362032 527054
rect 362268 526818 362352 527054
rect 362588 526818 362620 527054
rect 398000 527138 398032 527374
rect 398268 527138 398352 527374
rect 398588 527138 398620 527374
rect 398000 527054 398620 527138
rect 398000 526818 398032 527054
rect 398268 526818 398352 527054
rect 398588 526818 398620 527054
rect 434000 527138 434032 527374
rect 434268 527138 434352 527374
rect 434588 527138 434620 527374
rect 434000 527054 434620 527138
rect 434000 526818 434032 527054
rect 434268 526818 434352 527054
rect 434588 526818 434620 527054
rect 470000 527138 470032 527374
rect 470268 527138 470352 527374
rect 470588 527138 470620 527374
rect 470000 527054 470620 527138
rect 470000 526818 470032 527054
rect 470268 526818 470352 527054
rect 470588 526818 470620 527054
rect 506000 527138 506032 527374
rect 506268 527138 506352 527374
rect 506588 527138 506620 527374
rect 506000 527054 506620 527138
rect 506000 526818 506032 527054
rect 506268 526818 506352 527054
rect 506588 526818 506620 527054
rect 542000 527138 542032 527374
rect 542268 527138 542352 527374
rect 542588 527138 542620 527374
rect 542000 527054 542620 527138
rect 542000 526818 542032 527054
rect 542268 526818 542352 527054
rect 542588 526818 542620 527054
rect 571500 527138 571532 527374
rect 571768 527138 571852 527374
rect 572088 527138 572120 527374
rect 571500 527054 572120 527138
rect 571500 526818 571532 527054
rect 571768 526818 571852 527054
rect 572088 526818 572120 527054
rect -2006 523418 -1974 523654
rect -1738 523418 -1654 523654
rect -1418 523418 -1386 523654
rect -2006 523334 -1386 523418
rect -2006 523098 -1974 523334
rect -1738 523098 -1654 523334
rect -1418 523098 -1386 523334
rect 9084 523418 9116 523654
rect 9352 523418 9436 523654
rect 9672 523418 9704 523654
rect 9084 523334 9704 523418
rect 9084 523098 9116 523334
rect 9352 523098 9436 523334
rect 9672 523098 9704 523334
rect 56620 523418 56652 523654
rect 56888 523418 56972 523654
rect 57208 523418 57240 523654
rect 56620 523334 57240 523418
rect 56620 523098 56652 523334
rect 56888 523098 56972 523334
rect 57208 523098 57240 523334
rect 92620 523418 92652 523654
rect 92888 523418 92972 523654
rect 93208 523418 93240 523654
rect 92620 523334 93240 523418
rect 92620 523098 92652 523334
rect 92888 523098 92972 523334
rect 93208 523098 93240 523334
rect 128620 523418 128652 523654
rect 128888 523418 128972 523654
rect 129208 523418 129240 523654
rect 128620 523334 129240 523418
rect 128620 523098 128652 523334
rect 128888 523098 128972 523334
rect 129208 523098 129240 523334
rect 164620 523418 164652 523654
rect 164888 523418 164972 523654
rect 165208 523418 165240 523654
rect 164620 523334 165240 523418
rect 164620 523098 164652 523334
rect 164888 523098 164972 523334
rect 165208 523098 165240 523334
rect 200620 523418 200652 523654
rect 200888 523418 200972 523654
rect 201208 523418 201240 523654
rect 200620 523334 201240 523418
rect 200620 523098 200652 523334
rect 200888 523098 200972 523334
rect 201208 523098 201240 523334
rect 236620 523418 236652 523654
rect 236888 523418 236972 523654
rect 237208 523418 237240 523654
rect 236620 523334 237240 523418
rect 236620 523098 236652 523334
rect 236888 523098 236972 523334
rect 237208 523098 237240 523334
rect 272620 523418 272652 523654
rect 272888 523418 272972 523654
rect 273208 523418 273240 523654
rect 272620 523334 273240 523418
rect 272620 523098 272652 523334
rect 272888 523098 272972 523334
rect 273208 523098 273240 523334
rect 308620 523418 308652 523654
rect 308888 523418 308972 523654
rect 309208 523418 309240 523654
rect 308620 523334 309240 523418
rect 308620 523098 308652 523334
rect 308888 523098 308972 523334
rect 309208 523098 309240 523334
rect 344620 523418 344652 523654
rect 344888 523418 344972 523654
rect 345208 523418 345240 523654
rect 344620 523334 345240 523418
rect 344620 523098 344652 523334
rect 344888 523098 344972 523334
rect 345208 523098 345240 523334
rect 380620 523418 380652 523654
rect 380888 523418 380972 523654
rect 381208 523418 381240 523654
rect 380620 523334 381240 523418
rect 380620 523098 380652 523334
rect 380888 523098 380972 523334
rect 381208 523098 381240 523334
rect 416620 523418 416652 523654
rect 416888 523418 416972 523654
rect 417208 523418 417240 523654
rect 416620 523334 417240 523418
rect 416620 523098 416652 523334
rect 416888 523098 416972 523334
rect 417208 523098 417240 523334
rect 452620 523418 452652 523654
rect 452888 523418 452972 523654
rect 453208 523418 453240 523654
rect 452620 523334 453240 523418
rect 452620 523098 452652 523334
rect 452888 523098 452972 523334
rect 453208 523098 453240 523334
rect 488620 523418 488652 523654
rect 488888 523418 488972 523654
rect 489208 523418 489240 523654
rect 488620 523334 489240 523418
rect 488620 523098 488652 523334
rect 488888 523098 488972 523334
rect 489208 523098 489240 523334
rect 524620 523418 524652 523654
rect 524888 523418 524972 523654
rect 525208 523418 525240 523654
rect 524620 523334 525240 523418
rect 524620 523098 524652 523334
rect 524888 523098 524972 523334
rect 525208 523098 525240 523334
rect 560620 523418 560652 523654
rect 560888 523418 560972 523654
rect 561208 523418 561240 523654
rect 560620 523334 561240 523418
rect 560620 523098 560652 523334
rect 560888 523098 560972 523334
rect 561208 523098 561240 523334
rect 570260 523418 570292 523654
rect 570528 523418 570612 523654
rect 570848 523418 570880 523654
rect 570260 523334 570880 523418
rect 570260 523098 570292 523334
rect 570528 523098 570612 523334
rect 570848 523098 570880 523334
rect -2006 483654 -1386 523098
rect 580594 502254 581214 541698
rect 580594 502018 580626 502254
rect 580862 502018 580946 502254
rect 581182 502018 581214 502254
rect 580594 501934 581214 502018
rect 580594 501698 580626 501934
rect 580862 501698 580946 501934
rect 581182 501698 581214 501934
rect 60560 487374 60920 487406
rect 7844 487138 7876 487374
rect 8112 487138 8196 487374
rect 8432 487138 8464 487374
rect 7844 487054 8464 487138
rect 7844 486818 7876 487054
rect 8112 486818 8196 487054
rect 8432 486818 8464 487054
rect 38000 487138 38032 487374
rect 38268 487138 38352 487374
rect 38588 487138 38620 487374
rect 38000 487054 38620 487138
rect 38000 486818 38032 487054
rect 38268 486818 38352 487054
rect 38588 486818 38620 487054
rect 60560 487138 60622 487374
rect 60858 487138 60920 487374
rect 60560 487054 60920 487138
rect 60560 486818 60622 487054
rect 60858 486818 60920 487054
rect 60560 486786 60920 486818
rect 159036 487374 159396 487406
rect 185560 487374 185920 487406
rect 159036 487138 159098 487374
rect 159334 487138 159396 487374
rect 159036 487054 159396 487138
rect 159036 486818 159098 487054
rect 159334 486818 159396 487054
rect 182000 487138 182032 487374
rect 182268 487138 182352 487374
rect 182588 487138 182620 487374
rect 182000 487054 182620 487138
rect 182000 486818 182032 487054
rect 182268 486818 182352 487054
rect 182588 486818 182620 487054
rect 185560 487138 185622 487374
rect 185858 487138 185920 487374
rect 185560 487054 185920 487138
rect 185560 486818 185622 487054
rect 185858 486818 185920 487054
rect 159036 486786 159396 486818
rect 185560 486786 185920 486818
rect 284036 487374 284396 487406
rect 310560 487374 310920 487406
rect 284036 487138 284098 487374
rect 284334 487138 284396 487374
rect 284036 487054 284396 487138
rect 284036 486818 284098 487054
rect 284334 486818 284396 487054
rect 290000 487138 290032 487374
rect 290268 487138 290352 487374
rect 290588 487138 290620 487374
rect 290000 487054 290620 487138
rect 290000 486818 290032 487054
rect 290268 486818 290352 487054
rect 290588 486818 290620 487054
rect 310560 487138 310622 487374
rect 310858 487138 310920 487374
rect 310560 487054 310920 487138
rect 310560 486818 310622 487054
rect 310858 486818 310920 487054
rect 284036 486786 284396 486818
rect 310560 486786 310920 486818
rect 409036 487374 409396 487406
rect 436560 487374 436920 487406
rect 409036 487138 409098 487374
rect 409334 487138 409396 487374
rect 409036 487054 409396 487138
rect 409036 486818 409098 487054
rect 409334 486818 409396 487054
rect 434000 487138 434032 487374
rect 434268 487138 434352 487374
rect 434588 487138 434620 487374
rect 434000 487054 434620 487138
rect 434000 486818 434032 487054
rect 434268 486818 434352 487054
rect 434588 486818 434620 487054
rect 436560 487138 436622 487374
rect 436858 487138 436920 487374
rect 436560 487054 436920 487138
rect 436560 486818 436622 487054
rect 436858 486818 436920 487054
rect 409036 486786 409396 486818
rect 436560 486786 436920 486818
rect 535036 487374 535396 487406
rect 535036 487138 535098 487374
rect 535334 487138 535396 487374
rect 535036 487054 535396 487138
rect 535036 486818 535098 487054
rect 535334 486818 535396 487054
rect 542000 487138 542032 487374
rect 542268 487138 542352 487374
rect 542588 487138 542620 487374
rect 542000 487054 542620 487138
rect 542000 486818 542032 487054
rect 542268 486818 542352 487054
rect 542588 486818 542620 487054
rect 571500 487138 571532 487374
rect 571768 487138 571852 487374
rect 572088 487138 572120 487374
rect 571500 487054 572120 487138
rect 571500 486818 571532 487054
rect 571768 486818 571852 487054
rect 572088 486818 572120 487054
rect 535036 486786 535396 486818
rect 61280 483654 61640 483686
rect -2006 483418 -1974 483654
rect -1738 483418 -1654 483654
rect -1418 483418 -1386 483654
rect -2006 483334 -1386 483418
rect -2006 483098 -1974 483334
rect -1738 483098 -1654 483334
rect -1418 483098 -1386 483334
rect 9084 483418 9116 483654
rect 9352 483418 9436 483654
rect 9672 483418 9704 483654
rect 9084 483334 9704 483418
rect 9084 483098 9116 483334
rect 9352 483098 9436 483334
rect 9672 483098 9704 483334
rect 56620 483418 56652 483654
rect 56888 483418 56972 483654
rect 57208 483418 57240 483654
rect 56620 483334 57240 483418
rect 56620 483098 56652 483334
rect 56888 483098 56972 483334
rect 57208 483098 57240 483334
rect 61280 483418 61342 483654
rect 61578 483418 61640 483654
rect 61280 483334 61640 483418
rect 61280 483098 61342 483334
rect 61578 483098 61640 483334
rect -2006 443654 -1386 483098
rect 61280 483066 61640 483098
rect 158316 483654 158676 483686
rect 186280 483654 186640 483686
rect 158316 483418 158378 483654
rect 158614 483418 158676 483654
rect 158316 483334 158676 483418
rect 158316 483098 158378 483334
rect 158614 483098 158676 483334
rect 164620 483418 164652 483654
rect 164888 483418 164972 483654
rect 165208 483418 165240 483654
rect 164620 483334 165240 483418
rect 164620 483098 164652 483334
rect 164888 483098 164972 483334
rect 165208 483098 165240 483334
rect 186280 483418 186342 483654
rect 186578 483418 186640 483654
rect 186280 483334 186640 483418
rect 186280 483098 186342 483334
rect 186578 483098 186640 483334
rect 158316 483066 158676 483098
rect 186280 483066 186640 483098
rect 283316 483654 283676 483686
rect 311280 483654 311640 483686
rect 283316 483418 283378 483654
rect 283614 483418 283676 483654
rect 283316 483334 283676 483418
rect 283316 483098 283378 483334
rect 283614 483098 283676 483334
rect 308620 483418 308652 483654
rect 308888 483418 308972 483654
rect 309208 483418 309240 483654
rect 308620 483334 309240 483418
rect 308620 483098 308652 483334
rect 308888 483098 308972 483334
rect 309208 483098 309240 483334
rect 311280 483418 311342 483654
rect 311578 483418 311640 483654
rect 311280 483334 311640 483418
rect 311280 483098 311342 483334
rect 311578 483098 311640 483334
rect 283316 483066 283676 483098
rect 311280 483066 311640 483098
rect 408316 483654 408676 483686
rect 437280 483654 437640 483686
rect 408316 483418 408378 483654
rect 408614 483418 408676 483654
rect 408316 483334 408676 483418
rect 408316 483098 408378 483334
rect 408614 483098 408676 483334
rect 416620 483418 416652 483654
rect 416888 483418 416972 483654
rect 417208 483418 417240 483654
rect 416620 483334 417240 483418
rect 416620 483098 416652 483334
rect 416888 483098 416972 483334
rect 417208 483098 417240 483334
rect 437280 483418 437342 483654
rect 437578 483418 437640 483654
rect 437280 483334 437640 483418
rect 437280 483098 437342 483334
rect 437578 483098 437640 483334
rect 408316 483066 408676 483098
rect 437280 483066 437640 483098
rect 534316 483654 534676 483686
rect 534316 483418 534378 483654
rect 534614 483418 534676 483654
rect 534316 483334 534676 483418
rect 534316 483098 534378 483334
rect 534614 483098 534676 483334
rect 560620 483418 560652 483654
rect 560888 483418 560972 483654
rect 561208 483418 561240 483654
rect 560620 483334 561240 483418
rect 560620 483098 560652 483334
rect 560888 483098 560972 483334
rect 561208 483098 561240 483334
rect 570260 483418 570292 483654
rect 570528 483418 570612 483654
rect 570848 483418 570880 483654
rect 570260 483334 570880 483418
rect 570260 483098 570292 483334
rect 570528 483098 570612 483334
rect 570848 483098 570880 483334
rect 534316 483066 534676 483098
rect 580594 462254 581214 501698
rect 580594 462018 580626 462254
rect 580862 462018 580946 462254
rect 581182 462018 581214 462254
rect 580594 461934 581214 462018
rect 580594 461698 580626 461934
rect 580862 461698 580946 461934
rect 581182 461698 581214 461934
rect 60560 447374 60920 447406
rect 7844 447138 7876 447374
rect 8112 447138 8196 447374
rect 8432 447138 8464 447374
rect 7844 447054 8464 447138
rect 7844 446818 7876 447054
rect 8112 446818 8196 447054
rect 8432 446818 8464 447054
rect 38000 447138 38032 447374
rect 38268 447138 38352 447374
rect 38588 447138 38620 447374
rect 38000 447054 38620 447138
rect 38000 446818 38032 447054
rect 38268 446818 38352 447054
rect 38588 446818 38620 447054
rect 60560 447138 60622 447374
rect 60858 447138 60920 447374
rect 60560 447054 60920 447138
rect 60560 446818 60622 447054
rect 60858 446818 60920 447054
rect 60560 446786 60920 446818
rect 159036 447374 159396 447406
rect 185560 447374 185920 447406
rect 159036 447138 159098 447374
rect 159334 447138 159396 447374
rect 159036 447054 159396 447138
rect 159036 446818 159098 447054
rect 159334 446818 159396 447054
rect 182000 447138 182032 447374
rect 182268 447138 182352 447374
rect 182588 447138 182620 447374
rect 182000 447054 182620 447138
rect 182000 446818 182032 447054
rect 182268 446818 182352 447054
rect 182588 446818 182620 447054
rect 185560 447138 185622 447374
rect 185858 447138 185920 447374
rect 185560 447054 185920 447138
rect 185560 446818 185622 447054
rect 185858 446818 185920 447054
rect 159036 446786 159396 446818
rect 185560 446786 185920 446818
rect 284036 447374 284396 447406
rect 310560 447374 310920 447406
rect 284036 447138 284098 447374
rect 284334 447138 284396 447374
rect 284036 447054 284396 447138
rect 284036 446818 284098 447054
rect 284334 446818 284396 447054
rect 290000 447138 290032 447374
rect 290268 447138 290352 447374
rect 290588 447138 290620 447374
rect 290000 447054 290620 447138
rect 290000 446818 290032 447054
rect 290268 446818 290352 447054
rect 290588 446818 290620 447054
rect 310560 447138 310622 447374
rect 310858 447138 310920 447374
rect 310560 447054 310920 447138
rect 310560 446818 310622 447054
rect 310858 446818 310920 447054
rect 284036 446786 284396 446818
rect 310560 446786 310920 446818
rect 409036 447374 409396 447406
rect 436560 447374 436920 447406
rect 409036 447138 409098 447374
rect 409334 447138 409396 447374
rect 409036 447054 409396 447138
rect 409036 446818 409098 447054
rect 409334 446818 409396 447054
rect 434000 447138 434032 447374
rect 434268 447138 434352 447374
rect 434588 447138 434620 447374
rect 434000 447054 434620 447138
rect 434000 446818 434032 447054
rect 434268 446818 434352 447054
rect 434588 446818 434620 447054
rect 436560 447138 436622 447374
rect 436858 447138 436920 447374
rect 436560 447054 436920 447138
rect 436560 446818 436622 447054
rect 436858 446818 436920 447054
rect 409036 446786 409396 446818
rect 436560 446786 436920 446818
rect 535036 447374 535396 447406
rect 535036 447138 535098 447374
rect 535334 447138 535396 447374
rect 535036 447054 535396 447138
rect 535036 446818 535098 447054
rect 535334 446818 535396 447054
rect 542000 447138 542032 447374
rect 542268 447138 542352 447374
rect 542588 447138 542620 447374
rect 542000 447054 542620 447138
rect 542000 446818 542032 447054
rect 542268 446818 542352 447054
rect 542588 446818 542620 447054
rect 571500 447138 571532 447374
rect 571768 447138 571852 447374
rect 572088 447138 572120 447374
rect 571500 447054 572120 447138
rect 571500 446818 571532 447054
rect 571768 446818 571852 447054
rect 572088 446818 572120 447054
rect 535036 446786 535396 446818
rect 61280 443654 61640 443686
rect -2006 443418 -1974 443654
rect -1738 443418 -1654 443654
rect -1418 443418 -1386 443654
rect -2006 443334 -1386 443418
rect -2006 443098 -1974 443334
rect -1738 443098 -1654 443334
rect -1418 443098 -1386 443334
rect 9084 443418 9116 443654
rect 9352 443418 9436 443654
rect 9672 443418 9704 443654
rect 9084 443334 9704 443418
rect 9084 443098 9116 443334
rect 9352 443098 9436 443334
rect 9672 443098 9704 443334
rect 56620 443418 56652 443654
rect 56888 443418 56972 443654
rect 57208 443418 57240 443654
rect 56620 443334 57240 443418
rect 56620 443098 56652 443334
rect 56888 443098 56972 443334
rect 57208 443098 57240 443334
rect 61280 443418 61342 443654
rect 61578 443418 61640 443654
rect 61280 443334 61640 443418
rect 61280 443098 61342 443334
rect 61578 443098 61640 443334
rect -2006 403654 -1386 443098
rect 61280 443066 61640 443098
rect 158316 443654 158676 443686
rect 186280 443654 186640 443686
rect 158316 443418 158378 443654
rect 158614 443418 158676 443654
rect 158316 443334 158676 443418
rect 158316 443098 158378 443334
rect 158614 443098 158676 443334
rect 164620 443418 164652 443654
rect 164888 443418 164972 443654
rect 165208 443418 165240 443654
rect 164620 443334 165240 443418
rect 164620 443098 164652 443334
rect 164888 443098 164972 443334
rect 165208 443098 165240 443334
rect 186280 443418 186342 443654
rect 186578 443418 186640 443654
rect 186280 443334 186640 443418
rect 186280 443098 186342 443334
rect 186578 443098 186640 443334
rect 158316 443066 158676 443098
rect 186280 443066 186640 443098
rect 283316 443654 283676 443686
rect 311280 443654 311640 443686
rect 283316 443418 283378 443654
rect 283614 443418 283676 443654
rect 283316 443334 283676 443418
rect 283316 443098 283378 443334
rect 283614 443098 283676 443334
rect 308620 443418 308652 443654
rect 308888 443418 308972 443654
rect 309208 443418 309240 443654
rect 308620 443334 309240 443418
rect 308620 443098 308652 443334
rect 308888 443098 308972 443334
rect 309208 443098 309240 443334
rect 311280 443418 311342 443654
rect 311578 443418 311640 443654
rect 311280 443334 311640 443418
rect 311280 443098 311342 443334
rect 311578 443098 311640 443334
rect 283316 443066 283676 443098
rect 311280 443066 311640 443098
rect 408316 443654 408676 443686
rect 437280 443654 437640 443686
rect 408316 443418 408378 443654
rect 408614 443418 408676 443654
rect 408316 443334 408676 443418
rect 408316 443098 408378 443334
rect 408614 443098 408676 443334
rect 416620 443418 416652 443654
rect 416888 443418 416972 443654
rect 417208 443418 417240 443654
rect 416620 443334 417240 443418
rect 416620 443098 416652 443334
rect 416888 443098 416972 443334
rect 417208 443098 417240 443334
rect 437280 443418 437342 443654
rect 437578 443418 437640 443654
rect 437280 443334 437640 443418
rect 437280 443098 437342 443334
rect 437578 443098 437640 443334
rect 408316 443066 408676 443098
rect 437280 443066 437640 443098
rect 534316 443654 534676 443686
rect 534316 443418 534378 443654
rect 534614 443418 534676 443654
rect 534316 443334 534676 443418
rect 534316 443098 534378 443334
rect 534614 443098 534676 443334
rect 560620 443418 560652 443654
rect 560888 443418 560972 443654
rect 561208 443418 561240 443654
rect 560620 443334 561240 443418
rect 560620 443098 560652 443334
rect 560888 443098 560972 443334
rect 561208 443098 561240 443334
rect 570260 443418 570292 443654
rect 570528 443418 570612 443654
rect 570848 443418 570880 443654
rect 570260 443334 570880 443418
rect 570260 443098 570292 443334
rect 570528 443098 570612 443334
rect 570848 443098 570880 443334
rect 534316 443066 534676 443098
rect 61280 433244 61640 433300
rect 61280 433008 61342 433244
rect 61578 433008 61640 433244
rect 61280 432952 61640 433008
rect 62952 433244 63300 433300
rect 62952 433008 63008 433244
rect 63244 433008 63300 433244
rect 62952 432952 63300 433008
rect 281656 433244 282004 433300
rect 281656 433008 281712 433244
rect 281948 433008 282004 433244
rect 281656 432952 282004 433008
rect 283316 433244 283676 433300
rect 283316 433008 283378 433244
rect 283614 433008 283676 433244
rect 283316 432952 283676 433008
rect 311280 433244 311640 433300
rect 311280 433008 311342 433244
rect 311578 433008 311640 433244
rect 311280 432952 311640 433008
rect 312952 433244 313300 433300
rect 312952 433008 313008 433244
rect 313244 433008 313300 433244
rect 312952 432952 313300 433008
rect 532656 433244 533004 433300
rect 532656 433008 532712 433244
rect 532948 433008 533004 433244
rect 532656 432952 533004 433008
rect 534316 433244 534676 433300
rect 534316 433008 534378 433244
rect 534614 433008 534676 433244
rect 534316 432952 534676 433008
rect 157336 432564 157684 432620
rect 157336 432328 157392 432564
rect 157628 432328 157684 432564
rect 157336 432272 157684 432328
rect 159036 432564 159396 432620
rect 159036 432328 159098 432564
rect 159334 432328 159396 432564
rect 159036 432272 159396 432328
rect 185560 432564 185920 432620
rect 185560 432328 185622 432564
rect 185858 432328 185920 432564
rect 185560 432272 185920 432328
rect 187272 432564 187620 432620
rect 187272 432328 187328 432564
rect 187564 432328 187620 432564
rect 187272 432272 187620 432328
rect 407336 432564 407684 432620
rect 407336 432328 407392 432564
rect 407628 432328 407684 432564
rect 407336 432272 407684 432328
rect 409036 432564 409396 432620
rect 409036 432328 409098 432564
rect 409334 432328 409396 432564
rect 409036 432272 409396 432328
rect 436560 432564 436920 432620
rect 436560 432328 436622 432564
rect 436858 432328 436920 432564
rect 436560 432272 436920 432328
rect 438272 432564 438620 432620
rect 438272 432328 438328 432564
rect 438564 432328 438620 432564
rect 438272 432272 438620 432328
rect 580594 422254 581214 461698
rect 580594 422018 580626 422254
rect 580862 422018 580946 422254
rect 581182 422018 581214 422254
rect 580594 421934 581214 422018
rect 580594 421698 580626 421934
rect 580862 421698 580946 421934
rect 581182 421698 581214 421934
rect 7844 407138 7876 407374
rect 8112 407138 8196 407374
rect 8432 407138 8464 407374
rect 7844 407054 8464 407138
rect 7844 406818 7876 407054
rect 8112 406818 8196 407054
rect 8432 406818 8464 407054
rect 38000 407138 38032 407374
rect 38268 407138 38352 407374
rect 38588 407138 38620 407374
rect 38000 407054 38620 407138
rect 38000 406818 38032 407054
rect 38268 406818 38352 407054
rect 38588 406818 38620 407054
rect 74000 407138 74032 407374
rect 74268 407138 74352 407374
rect 74588 407138 74620 407374
rect 74000 407054 74620 407138
rect 74000 406818 74032 407054
rect 74268 406818 74352 407054
rect 74588 406818 74620 407054
rect 110000 407138 110032 407374
rect 110268 407138 110352 407374
rect 110588 407138 110620 407374
rect 110000 407054 110620 407138
rect 110000 406818 110032 407054
rect 110268 406818 110352 407054
rect 110588 406818 110620 407054
rect 146000 407138 146032 407374
rect 146268 407138 146352 407374
rect 146588 407138 146620 407374
rect 146000 407054 146620 407138
rect 146000 406818 146032 407054
rect 146268 406818 146352 407054
rect 146588 406818 146620 407054
rect 182000 407138 182032 407374
rect 182268 407138 182352 407374
rect 182588 407138 182620 407374
rect 182000 407054 182620 407138
rect 182000 406818 182032 407054
rect 182268 406818 182352 407054
rect 182588 406818 182620 407054
rect 218000 407138 218032 407374
rect 218268 407138 218352 407374
rect 218588 407138 218620 407374
rect 218000 407054 218620 407138
rect 218000 406818 218032 407054
rect 218268 406818 218352 407054
rect 218588 406818 218620 407054
rect 254000 407138 254032 407374
rect 254268 407138 254352 407374
rect 254588 407138 254620 407374
rect 254000 407054 254620 407138
rect 254000 406818 254032 407054
rect 254268 406818 254352 407054
rect 254588 406818 254620 407054
rect 290000 407138 290032 407374
rect 290268 407138 290352 407374
rect 290588 407138 290620 407374
rect 290000 407054 290620 407138
rect 290000 406818 290032 407054
rect 290268 406818 290352 407054
rect 290588 406818 290620 407054
rect 326000 407138 326032 407374
rect 326268 407138 326352 407374
rect 326588 407138 326620 407374
rect 326000 407054 326620 407138
rect 326000 406818 326032 407054
rect 326268 406818 326352 407054
rect 326588 406818 326620 407054
rect 362000 407138 362032 407374
rect 362268 407138 362352 407374
rect 362588 407138 362620 407374
rect 362000 407054 362620 407138
rect 362000 406818 362032 407054
rect 362268 406818 362352 407054
rect 362588 406818 362620 407054
rect 398000 407138 398032 407374
rect 398268 407138 398352 407374
rect 398588 407138 398620 407374
rect 398000 407054 398620 407138
rect 398000 406818 398032 407054
rect 398268 406818 398352 407054
rect 398588 406818 398620 407054
rect 434000 407138 434032 407374
rect 434268 407138 434352 407374
rect 434588 407138 434620 407374
rect 434000 407054 434620 407138
rect 434000 406818 434032 407054
rect 434268 406818 434352 407054
rect 434588 406818 434620 407054
rect 470000 407138 470032 407374
rect 470268 407138 470352 407374
rect 470588 407138 470620 407374
rect 470000 407054 470620 407138
rect 470000 406818 470032 407054
rect 470268 406818 470352 407054
rect 470588 406818 470620 407054
rect 506000 407138 506032 407374
rect 506268 407138 506352 407374
rect 506588 407138 506620 407374
rect 506000 407054 506620 407138
rect 506000 406818 506032 407054
rect 506268 406818 506352 407054
rect 506588 406818 506620 407054
rect 542000 407138 542032 407374
rect 542268 407138 542352 407374
rect 542588 407138 542620 407374
rect 542000 407054 542620 407138
rect 542000 406818 542032 407054
rect 542268 406818 542352 407054
rect 542588 406818 542620 407054
rect 571500 407138 571532 407374
rect 571768 407138 571852 407374
rect 572088 407138 572120 407374
rect 571500 407054 572120 407138
rect 571500 406818 571532 407054
rect 571768 406818 571852 407054
rect 572088 406818 572120 407054
rect -2006 403418 -1974 403654
rect -1738 403418 -1654 403654
rect -1418 403418 -1386 403654
rect -2006 403334 -1386 403418
rect -2006 403098 -1974 403334
rect -1738 403098 -1654 403334
rect -1418 403098 -1386 403334
rect 9084 403418 9116 403654
rect 9352 403418 9436 403654
rect 9672 403418 9704 403654
rect 9084 403334 9704 403418
rect 9084 403098 9116 403334
rect 9352 403098 9436 403334
rect 9672 403098 9704 403334
rect 56620 403418 56652 403654
rect 56888 403418 56972 403654
rect 57208 403418 57240 403654
rect 56620 403334 57240 403418
rect 56620 403098 56652 403334
rect 56888 403098 56972 403334
rect 57208 403098 57240 403334
rect 92620 403418 92652 403654
rect 92888 403418 92972 403654
rect 93208 403418 93240 403654
rect 92620 403334 93240 403418
rect 92620 403098 92652 403334
rect 92888 403098 92972 403334
rect 93208 403098 93240 403334
rect 128620 403418 128652 403654
rect 128888 403418 128972 403654
rect 129208 403418 129240 403654
rect 128620 403334 129240 403418
rect 128620 403098 128652 403334
rect 128888 403098 128972 403334
rect 129208 403098 129240 403334
rect 164620 403418 164652 403654
rect 164888 403418 164972 403654
rect 165208 403418 165240 403654
rect 164620 403334 165240 403418
rect 164620 403098 164652 403334
rect 164888 403098 164972 403334
rect 165208 403098 165240 403334
rect 200620 403418 200652 403654
rect 200888 403418 200972 403654
rect 201208 403418 201240 403654
rect 200620 403334 201240 403418
rect 200620 403098 200652 403334
rect 200888 403098 200972 403334
rect 201208 403098 201240 403334
rect 236620 403418 236652 403654
rect 236888 403418 236972 403654
rect 237208 403418 237240 403654
rect 236620 403334 237240 403418
rect 236620 403098 236652 403334
rect 236888 403098 236972 403334
rect 237208 403098 237240 403334
rect 272620 403418 272652 403654
rect 272888 403418 272972 403654
rect 273208 403418 273240 403654
rect 272620 403334 273240 403418
rect 272620 403098 272652 403334
rect 272888 403098 272972 403334
rect 273208 403098 273240 403334
rect 308620 403418 308652 403654
rect 308888 403418 308972 403654
rect 309208 403418 309240 403654
rect 308620 403334 309240 403418
rect 308620 403098 308652 403334
rect 308888 403098 308972 403334
rect 309208 403098 309240 403334
rect 344620 403418 344652 403654
rect 344888 403418 344972 403654
rect 345208 403418 345240 403654
rect 344620 403334 345240 403418
rect 344620 403098 344652 403334
rect 344888 403098 344972 403334
rect 345208 403098 345240 403334
rect 380620 403418 380652 403654
rect 380888 403418 380972 403654
rect 381208 403418 381240 403654
rect 380620 403334 381240 403418
rect 380620 403098 380652 403334
rect 380888 403098 380972 403334
rect 381208 403098 381240 403334
rect 416620 403418 416652 403654
rect 416888 403418 416972 403654
rect 417208 403418 417240 403654
rect 416620 403334 417240 403418
rect 416620 403098 416652 403334
rect 416888 403098 416972 403334
rect 417208 403098 417240 403334
rect 452620 403418 452652 403654
rect 452888 403418 452972 403654
rect 453208 403418 453240 403654
rect 452620 403334 453240 403418
rect 452620 403098 452652 403334
rect 452888 403098 452972 403334
rect 453208 403098 453240 403334
rect 488620 403418 488652 403654
rect 488888 403418 488972 403654
rect 489208 403418 489240 403654
rect 488620 403334 489240 403418
rect 488620 403098 488652 403334
rect 488888 403098 488972 403334
rect 489208 403098 489240 403334
rect 524620 403418 524652 403654
rect 524888 403418 524972 403654
rect 525208 403418 525240 403654
rect 524620 403334 525240 403418
rect 524620 403098 524652 403334
rect 524888 403098 524972 403334
rect 525208 403098 525240 403334
rect 560620 403418 560652 403654
rect 560888 403418 560972 403654
rect 561208 403418 561240 403654
rect 560620 403334 561240 403418
rect 560620 403098 560652 403334
rect 560888 403098 560972 403334
rect 561208 403098 561240 403334
rect 570260 403418 570292 403654
rect 570528 403418 570612 403654
rect 570848 403418 570880 403654
rect 570260 403334 570880 403418
rect 570260 403098 570292 403334
rect 570528 403098 570612 403334
rect 570848 403098 570880 403334
rect -2006 363654 -1386 403098
rect 580594 382254 581214 421698
rect 580594 382018 580626 382254
rect 580862 382018 580946 382254
rect 581182 382018 581214 382254
rect 580594 381934 581214 382018
rect 580594 381698 580626 381934
rect 580862 381698 580946 381934
rect 581182 381698 581214 381934
rect 7844 367138 7876 367374
rect 8112 367138 8196 367374
rect 8432 367138 8464 367374
rect 7844 367054 8464 367138
rect 7844 366818 7876 367054
rect 8112 366818 8196 367054
rect 8432 366818 8464 367054
rect 38000 367138 38032 367374
rect 38268 367138 38352 367374
rect 38588 367138 38620 367374
rect 38000 367054 38620 367138
rect 38000 366818 38032 367054
rect 38268 366818 38352 367054
rect 38588 366818 38620 367054
rect 74000 367138 74032 367374
rect 74268 367138 74352 367374
rect 74588 367138 74620 367374
rect 74000 367054 74620 367138
rect 74000 366818 74032 367054
rect 74268 366818 74352 367054
rect 74588 366818 74620 367054
rect 110000 367138 110032 367374
rect 110268 367138 110352 367374
rect 110588 367138 110620 367374
rect 110000 367054 110620 367138
rect 110000 366818 110032 367054
rect 110268 366818 110352 367054
rect 110588 366818 110620 367054
rect 146000 367138 146032 367374
rect 146268 367138 146352 367374
rect 146588 367138 146620 367374
rect 146000 367054 146620 367138
rect 146000 366818 146032 367054
rect 146268 366818 146352 367054
rect 146588 366818 146620 367054
rect 182000 367138 182032 367374
rect 182268 367138 182352 367374
rect 182588 367138 182620 367374
rect 182000 367054 182620 367138
rect 182000 366818 182032 367054
rect 182268 366818 182352 367054
rect 182588 366818 182620 367054
rect 218000 367138 218032 367374
rect 218268 367138 218352 367374
rect 218588 367138 218620 367374
rect 218000 367054 218620 367138
rect 218000 366818 218032 367054
rect 218268 366818 218352 367054
rect 218588 366818 218620 367054
rect 254000 367138 254032 367374
rect 254268 367138 254352 367374
rect 254588 367138 254620 367374
rect 254000 367054 254620 367138
rect 254000 366818 254032 367054
rect 254268 366818 254352 367054
rect 254588 366818 254620 367054
rect 290000 367138 290032 367374
rect 290268 367138 290352 367374
rect 290588 367138 290620 367374
rect 290000 367054 290620 367138
rect 290000 366818 290032 367054
rect 290268 366818 290352 367054
rect 290588 366818 290620 367054
rect 326000 367138 326032 367374
rect 326268 367138 326352 367374
rect 326588 367138 326620 367374
rect 326000 367054 326620 367138
rect 326000 366818 326032 367054
rect 326268 366818 326352 367054
rect 326588 366818 326620 367054
rect 362000 367138 362032 367374
rect 362268 367138 362352 367374
rect 362588 367138 362620 367374
rect 362000 367054 362620 367138
rect 362000 366818 362032 367054
rect 362268 366818 362352 367054
rect 362588 366818 362620 367054
rect 398000 367138 398032 367374
rect 398268 367138 398352 367374
rect 398588 367138 398620 367374
rect 398000 367054 398620 367138
rect 398000 366818 398032 367054
rect 398268 366818 398352 367054
rect 398588 366818 398620 367054
rect 434000 367138 434032 367374
rect 434268 367138 434352 367374
rect 434588 367138 434620 367374
rect 434000 367054 434620 367138
rect 434000 366818 434032 367054
rect 434268 366818 434352 367054
rect 434588 366818 434620 367054
rect 470000 367138 470032 367374
rect 470268 367138 470352 367374
rect 470588 367138 470620 367374
rect 470000 367054 470620 367138
rect 470000 366818 470032 367054
rect 470268 366818 470352 367054
rect 470588 366818 470620 367054
rect 506000 367138 506032 367374
rect 506268 367138 506352 367374
rect 506588 367138 506620 367374
rect 506000 367054 506620 367138
rect 506000 366818 506032 367054
rect 506268 366818 506352 367054
rect 506588 366818 506620 367054
rect 542000 367138 542032 367374
rect 542268 367138 542352 367374
rect 542588 367138 542620 367374
rect 542000 367054 542620 367138
rect 542000 366818 542032 367054
rect 542268 366818 542352 367054
rect 542588 366818 542620 367054
rect 571500 367138 571532 367374
rect 571768 367138 571852 367374
rect 572088 367138 572120 367374
rect 571500 367054 572120 367138
rect 571500 366818 571532 367054
rect 571768 366818 571852 367054
rect 572088 366818 572120 367054
rect -2006 363418 -1974 363654
rect -1738 363418 -1654 363654
rect -1418 363418 -1386 363654
rect -2006 363334 -1386 363418
rect -2006 363098 -1974 363334
rect -1738 363098 -1654 363334
rect -1418 363098 -1386 363334
rect 9084 363418 9116 363654
rect 9352 363418 9436 363654
rect 9672 363418 9704 363654
rect 9084 363334 9704 363418
rect 9084 363098 9116 363334
rect 9352 363098 9436 363334
rect 9672 363098 9704 363334
rect 56620 363418 56652 363654
rect 56888 363418 56972 363654
rect 57208 363418 57240 363654
rect 56620 363334 57240 363418
rect 56620 363098 56652 363334
rect 56888 363098 56972 363334
rect 57208 363098 57240 363334
rect 92620 363418 92652 363654
rect 92888 363418 92972 363654
rect 93208 363418 93240 363654
rect 92620 363334 93240 363418
rect 92620 363098 92652 363334
rect 92888 363098 92972 363334
rect 93208 363098 93240 363334
rect 128620 363418 128652 363654
rect 128888 363418 128972 363654
rect 129208 363418 129240 363654
rect 128620 363334 129240 363418
rect 128620 363098 128652 363334
rect 128888 363098 128972 363334
rect 129208 363098 129240 363334
rect 164620 363418 164652 363654
rect 164888 363418 164972 363654
rect 165208 363418 165240 363654
rect 164620 363334 165240 363418
rect 164620 363098 164652 363334
rect 164888 363098 164972 363334
rect 165208 363098 165240 363334
rect 200620 363418 200652 363654
rect 200888 363418 200972 363654
rect 201208 363418 201240 363654
rect 200620 363334 201240 363418
rect 200620 363098 200652 363334
rect 200888 363098 200972 363334
rect 201208 363098 201240 363334
rect 236620 363418 236652 363654
rect 236888 363418 236972 363654
rect 237208 363418 237240 363654
rect 236620 363334 237240 363418
rect 236620 363098 236652 363334
rect 236888 363098 236972 363334
rect 237208 363098 237240 363334
rect 272620 363418 272652 363654
rect 272888 363418 272972 363654
rect 273208 363418 273240 363654
rect 272620 363334 273240 363418
rect 272620 363098 272652 363334
rect 272888 363098 272972 363334
rect 273208 363098 273240 363334
rect 308620 363418 308652 363654
rect 308888 363418 308972 363654
rect 309208 363418 309240 363654
rect 308620 363334 309240 363418
rect 308620 363098 308652 363334
rect 308888 363098 308972 363334
rect 309208 363098 309240 363334
rect 344620 363418 344652 363654
rect 344888 363418 344972 363654
rect 345208 363418 345240 363654
rect 344620 363334 345240 363418
rect 344620 363098 344652 363334
rect 344888 363098 344972 363334
rect 345208 363098 345240 363334
rect 380620 363418 380652 363654
rect 380888 363418 380972 363654
rect 381208 363418 381240 363654
rect 380620 363334 381240 363418
rect 380620 363098 380652 363334
rect 380888 363098 380972 363334
rect 381208 363098 381240 363334
rect 416620 363418 416652 363654
rect 416888 363418 416972 363654
rect 417208 363418 417240 363654
rect 416620 363334 417240 363418
rect 416620 363098 416652 363334
rect 416888 363098 416972 363334
rect 417208 363098 417240 363334
rect 452620 363418 452652 363654
rect 452888 363418 452972 363654
rect 453208 363418 453240 363654
rect 452620 363334 453240 363418
rect 452620 363098 452652 363334
rect 452888 363098 452972 363334
rect 453208 363098 453240 363334
rect 488620 363418 488652 363654
rect 488888 363418 488972 363654
rect 489208 363418 489240 363654
rect 488620 363334 489240 363418
rect 488620 363098 488652 363334
rect 488888 363098 488972 363334
rect 489208 363098 489240 363334
rect 524620 363418 524652 363654
rect 524888 363418 524972 363654
rect 525208 363418 525240 363654
rect 524620 363334 525240 363418
rect 524620 363098 524652 363334
rect 524888 363098 524972 363334
rect 525208 363098 525240 363334
rect 560620 363418 560652 363654
rect 560888 363418 560972 363654
rect 561208 363418 561240 363654
rect 560620 363334 561240 363418
rect 560620 363098 560652 363334
rect 560888 363098 560972 363334
rect 561208 363098 561240 363334
rect 570260 363418 570292 363654
rect 570528 363418 570612 363654
rect 570848 363418 570880 363654
rect 570260 363334 570880 363418
rect 570260 363098 570292 363334
rect 570528 363098 570612 363334
rect 570848 363098 570880 363334
rect -2006 323654 -1386 363098
rect 580594 342254 581214 381698
rect 580594 342018 580626 342254
rect 580862 342018 580946 342254
rect 581182 342018 581214 342254
rect 580594 341934 581214 342018
rect 580594 341698 580626 341934
rect 580862 341698 580946 341934
rect 581182 341698 581214 341934
rect 7844 327138 7876 327374
rect 8112 327138 8196 327374
rect 8432 327138 8464 327374
rect 7844 327054 8464 327138
rect 7844 326818 7876 327054
rect 8112 326818 8196 327054
rect 8432 326818 8464 327054
rect 38000 327138 38032 327374
rect 38268 327138 38352 327374
rect 38588 327138 38620 327374
rect 38000 327054 38620 327138
rect 38000 326818 38032 327054
rect 38268 326818 38352 327054
rect 38588 326818 38620 327054
rect 74000 327138 74032 327374
rect 74268 327138 74352 327374
rect 74588 327138 74620 327374
rect 74000 327054 74620 327138
rect 74000 326818 74032 327054
rect 74268 326818 74352 327054
rect 74588 326818 74620 327054
rect 110000 327138 110032 327374
rect 110268 327138 110352 327374
rect 110588 327138 110620 327374
rect 110000 327054 110620 327138
rect 110000 326818 110032 327054
rect 110268 326818 110352 327054
rect 110588 326818 110620 327054
rect 146000 327138 146032 327374
rect 146268 327138 146352 327374
rect 146588 327138 146620 327374
rect 146000 327054 146620 327138
rect 146000 326818 146032 327054
rect 146268 326818 146352 327054
rect 146588 326818 146620 327054
rect 182000 327138 182032 327374
rect 182268 327138 182352 327374
rect 182588 327138 182620 327374
rect 182000 327054 182620 327138
rect 182000 326818 182032 327054
rect 182268 326818 182352 327054
rect 182588 326818 182620 327054
rect 218000 327138 218032 327374
rect 218268 327138 218352 327374
rect 218588 327138 218620 327374
rect 218000 327054 218620 327138
rect 218000 326818 218032 327054
rect 218268 326818 218352 327054
rect 218588 326818 218620 327054
rect 254000 327138 254032 327374
rect 254268 327138 254352 327374
rect 254588 327138 254620 327374
rect 254000 327054 254620 327138
rect 254000 326818 254032 327054
rect 254268 326818 254352 327054
rect 254588 326818 254620 327054
rect 290000 327138 290032 327374
rect 290268 327138 290352 327374
rect 290588 327138 290620 327374
rect 290000 327054 290620 327138
rect 290000 326818 290032 327054
rect 290268 326818 290352 327054
rect 290588 326818 290620 327054
rect 326000 327138 326032 327374
rect 326268 327138 326352 327374
rect 326588 327138 326620 327374
rect 326000 327054 326620 327138
rect 326000 326818 326032 327054
rect 326268 326818 326352 327054
rect 326588 326818 326620 327054
rect 362000 327138 362032 327374
rect 362268 327138 362352 327374
rect 362588 327138 362620 327374
rect 362000 327054 362620 327138
rect 362000 326818 362032 327054
rect 362268 326818 362352 327054
rect 362588 326818 362620 327054
rect 398000 327138 398032 327374
rect 398268 327138 398352 327374
rect 398588 327138 398620 327374
rect 398000 327054 398620 327138
rect 398000 326818 398032 327054
rect 398268 326818 398352 327054
rect 398588 326818 398620 327054
rect 434000 327138 434032 327374
rect 434268 327138 434352 327374
rect 434588 327138 434620 327374
rect 434000 327054 434620 327138
rect 434000 326818 434032 327054
rect 434268 326818 434352 327054
rect 434588 326818 434620 327054
rect 470000 327138 470032 327374
rect 470268 327138 470352 327374
rect 470588 327138 470620 327374
rect 470000 327054 470620 327138
rect 470000 326818 470032 327054
rect 470268 326818 470352 327054
rect 470588 326818 470620 327054
rect 506000 327138 506032 327374
rect 506268 327138 506352 327374
rect 506588 327138 506620 327374
rect 506000 327054 506620 327138
rect 506000 326818 506032 327054
rect 506268 326818 506352 327054
rect 506588 326818 506620 327054
rect 542000 327138 542032 327374
rect 542268 327138 542352 327374
rect 542588 327138 542620 327374
rect 542000 327054 542620 327138
rect 542000 326818 542032 327054
rect 542268 326818 542352 327054
rect 542588 326818 542620 327054
rect 571500 327138 571532 327374
rect 571768 327138 571852 327374
rect 572088 327138 572120 327374
rect 571500 327054 572120 327138
rect 571500 326818 571532 327054
rect 571768 326818 571852 327054
rect 572088 326818 572120 327054
rect -2006 323418 -1974 323654
rect -1738 323418 -1654 323654
rect -1418 323418 -1386 323654
rect -2006 323334 -1386 323418
rect -2006 323098 -1974 323334
rect -1738 323098 -1654 323334
rect -1418 323098 -1386 323334
rect 9084 323418 9116 323654
rect 9352 323418 9436 323654
rect 9672 323418 9704 323654
rect 9084 323334 9704 323418
rect 9084 323098 9116 323334
rect 9352 323098 9436 323334
rect 9672 323098 9704 323334
rect 56620 323418 56652 323654
rect 56888 323418 56972 323654
rect 57208 323418 57240 323654
rect 56620 323334 57240 323418
rect 56620 323098 56652 323334
rect 56888 323098 56972 323334
rect 57208 323098 57240 323334
rect 92620 323418 92652 323654
rect 92888 323418 92972 323654
rect 93208 323418 93240 323654
rect 92620 323334 93240 323418
rect 92620 323098 92652 323334
rect 92888 323098 92972 323334
rect 93208 323098 93240 323334
rect 128620 323418 128652 323654
rect 128888 323418 128972 323654
rect 129208 323418 129240 323654
rect 128620 323334 129240 323418
rect 128620 323098 128652 323334
rect 128888 323098 128972 323334
rect 129208 323098 129240 323334
rect 164620 323418 164652 323654
rect 164888 323418 164972 323654
rect 165208 323418 165240 323654
rect 164620 323334 165240 323418
rect 164620 323098 164652 323334
rect 164888 323098 164972 323334
rect 165208 323098 165240 323334
rect 200620 323418 200652 323654
rect 200888 323418 200972 323654
rect 201208 323418 201240 323654
rect 200620 323334 201240 323418
rect 200620 323098 200652 323334
rect 200888 323098 200972 323334
rect 201208 323098 201240 323334
rect 236620 323418 236652 323654
rect 236888 323418 236972 323654
rect 237208 323418 237240 323654
rect 236620 323334 237240 323418
rect 236620 323098 236652 323334
rect 236888 323098 236972 323334
rect 237208 323098 237240 323334
rect 272620 323418 272652 323654
rect 272888 323418 272972 323654
rect 273208 323418 273240 323654
rect 272620 323334 273240 323418
rect 272620 323098 272652 323334
rect 272888 323098 272972 323334
rect 273208 323098 273240 323334
rect 308620 323418 308652 323654
rect 308888 323418 308972 323654
rect 309208 323418 309240 323654
rect 308620 323334 309240 323418
rect 308620 323098 308652 323334
rect 308888 323098 308972 323334
rect 309208 323098 309240 323334
rect 344620 323418 344652 323654
rect 344888 323418 344972 323654
rect 345208 323418 345240 323654
rect 344620 323334 345240 323418
rect 344620 323098 344652 323334
rect 344888 323098 344972 323334
rect 345208 323098 345240 323334
rect 380620 323418 380652 323654
rect 380888 323418 380972 323654
rect 381208 323418 381240 323654
rect 380620 323334 381240 323418
rect 380620 323098 380652 323334
rect 380888 323098 380972 323334
rect 381208 323098 381240 323334
rect 416620 323418 416652 323654
rect 416888 323418 416972 323654
rect 417208 323418 417240 323654
rect 416620 323334 417240 323418
rect 416620 323098 416652 323334
rect 416888 323098 416972 323334
rect 417208 323098 417240 323334
rect 452620 323418 452652 323654
rect 452888 323418 452972 323654
rect 453208 323418 453240 323654
rect 452620 323334 453240 323418
rect 452620 323098 452652 323334
rect 452888 323098 452972 323334
rect 453208 323098 453240 323334
rect 488620 323418 488652 323654
rect 488888 323418 488972 323654
rect 489208 323418 489240 323654
rect 488620 323334 489240 323418
rect 488620 323098 488652 323334
rect 488888 323098 488972 323334
rect 489208 323098 489240 323334
rect 524620 323418 524652 323654
rect 524888 323418 524972 323654
rect 525208 323418 525240 323654
rect 524620 323334 525240 323418
rect 524620 323098 524652 323334
rect 524888 323098 524972 323334
rect 525208 323098 525240 323334
rect 560620 323418 560652 323654
rect 560888 323418 560972 323654
rect 561208 323418 561240 323654
rect 560620 323334 561240 323418
rect 560620 323098 560652 323334
rect 560888 323098 560972 323334
rect 561208 323098 561240 323334
rect 570260 323418 570292 323654
rect 570528 323418 570612 323654
rect 570848 323418 570880 323654
rect 570260 323334 570880 323418
rect 570260 323098 570292 323334
rect 570528 323098 570612 323334
rect 570848 323098 570880 323334
rect -2006 283654 -1386 323098
rect 580594 302254 581214 341698
rect 580594 302018 580626 302254
rect 580862 302018 580946 302254
rect 581182 302018 581214 302254
rect 580594 301934 581214 302018
rect 580594 301698 580626 301934
rect 580862 301698 580946 301934
rect 581182 301698 581214 301934
rect 7844 287138 7876 287374
rect 8112 287138 8196 287374
rect 8432 287138 8464 287374
rect 7844 287054 8464 287138
rect 7844 286818 7876 287054
rect 8112 286818 8196 287054
rect 8432 286818 8464 287054
rect 38000 287138 38032 287374
rect 38268 287138 38352 287374
rect 38588 287138 38620 287374
rect 38000 287054 38620 287138
rect 38000 286818 38032 287054
rect 38268 286818 38352 287054
rect 38588 286818 38620 287054
rect 74000 287138 74032 287374
rect 74268 287138 74352 287374
rect 74588 287138 74620 287374
rect 74000 287054 74620 287138
rect 74000 286818 74032 287054
rect 74268 286818 74352 287054
rect 74588 286818 74620 287054
rect 110000 287138 110032 287374
rect 110268 287138 110352 287374
rect 110588 287138 110620 287374
rect 110000 287054 110620 287138
rect 110000 286818 110032 287054
rect 110268 286818 110352 287054
rect 110588 286818 110620 287054
rect 146000 287138 146032 287374
rect 146268 287138 146352 287374
rect 146588 287138 146620 287374
rect 146000 287054 146620 287138
rect 146000 286818 146032 287054
rect 146268 286818 146352 287054
rect 146588 286818 146620 287054
rect 182000 287138 182032 287374
rect 182268 287138 182352 287374
rect 182588 287138 182620 287374
rect 182000 287054 182620 287138
rect 182000 286818 182032 287054
rect 182268 286818 182352 287054
rect 182588 286818 182620 287054
rect 218000 287138 218032 287374
rect 218268 287138 218352 287374
rect 218588 287138 218620 287374
rect 218000 287054 218620 287138
rect 218000 286818 218032 287054
rect 218268 286818 218352 287054
rect 218588 286818 218620 287054
rect 254000 287138 254032 287374
rect 254268 287138 254352 287374
rect 254588 287138 254620 287374
rect 254000 287054 254620 287138
rect 254000 286818 254032 287054
rect 254268 286818 254352 287054
rect 254588 286818 254620 287054
rect 290000 287138 290032 287374
rect 290268 287138 290352 287374
rect 290588 287138 290620 287374
rect 290000 287054 290620 287138
rect 290000 286818 290032 287054
rect 290268 286818 290352 287054
rect 290588 286818 290620 287054
rect 326000 287138 326032 287374
rect 326268 287138 326352 287374
rect 326588 287138 326620 287374
rect 326000 287054 326620 287138
rect 326000 286818 326032 287054
rect 326268 286818 326352 287054
rect 326588 286818 326620 287054
rect 362000 287138 362032 287374
rect 362268 287138 362352 287374
rect 362588 287138 362620 287374
rect 362000 287054 362620 287138
rect 362000 286818 362032 287054
rect 362268 286818 362352 287054
rect 362588 286818 362620 287054
rect 398000 287138 398032 287374
rect 398268 287138 398352 287374
rect 398588 287138 398620 287374
rect 398000 287054 398620 287138
rect 398000 286818 398032 287054
rect 398268 286818 398352 287054
rect 398588 286818 398620 287054
rect 434000 287138 434032 287374
rect 434268 287138 434352 287374
rect 434588 287138 434620 287374
rect 434000 287054 434620 287138
rect 434000 286818 434032 287054
rect 434268 286818 434352 287054
rect 434588 286818 434620 287054
rect 470000 287138 470032 287374
rect 470268 287138 470352 287374
rect 470588 287138 470620 287374
rect 470000 287054 470620 287138
rect 470000 286818 470032 287054
rect 470268 286818 470352 287054
rect 470588 286818 470620 287054
rect 506000 287138 506032 287374
rect 506268 287138 506352 287374
rect 506588 287138 506620 287374
rect 506000 287054 506620 287138
rect 506000 286818 506032 287054
rect 506268 286818 506352 287054
rect 506588 286818 506620 287054
rect 542000 287138 542032 287374
rect 542268 287138 542352 287374
rect 542588 287138 542620 287374
rect 542000 287054 542620 287138
rect 542000 286818 542032 287054
rect 542268 286818 542352 287054
rect 542588 286818 542620 287054
rect 571500 287138 571532 287374
rect 571768 287138 571852 287374
rect 572088 287138 572120 287374
rect 571500 287054 572120 287138
rect 571500 286818 571532 287054
rect 571768 286818 571852 287054
rect 572088 286818 572120 287054
rect -2006 283418 -1974 283654
rect -1738 283418 -1654 283654
rect -1418 283418 -1386 283654
rect -2006 283334 -1386 283418
rect -2006 283098 -1974 283334
rect -1738 283098 -1654 283334
rect -1418 283098 -1386 283334
rect 9084 283418 9116 283654
rect 9352 283418 9436 283654
rect 9672 283418 9704 283654
rect 9084 283334 9704 283418
rect 9084 283098 9116 283334
rect 9352 283098 9436 283334
rect 9672 283098 9704 283334
rect 56620 283418 56652 283654
rect 56888 283418 56972 283654
rect 57208 283418 57240 283654
rect 56620 283334 57240 283418
rect 56620 283098 56652 283334
rect 56888 283098 56972 283334
rect 57208 283098 57240 283334
rect 92620 283418 92652 283654
rect 92888 283418 92972 283654
rect 93208 283418 93240 283654
rect 92620 283334 93240 283418
rect 92620 283098 92652 283334
rect 92888 283098 92972 283334
rect 93208 283098 93240 283334
rect 128620 283418 128652 283654
rect 128888 283418 128972 283654
rect 129208 283418 129240 283654
rect 128620 283334 129240 283418
rect 128620 283098 128652 283334
rect 128888 283098 128972 283334
rect 129208 283098 129240 283334
rect 164620 283418 164652 283654
rect 164888 283418 164972 283654
rect 165208 283418 165240 283654
rect 164620 283334 165240 283418
rect 164620 283098 164652 283334
rect 164888 283098 164972 283334
rect 165208 283098 165240 283334
rect 200620 283418 200652 283654
rect 200888 283418 200972 283654
rect 201208 283418 201240 283654
rect 200620 283334 201240 283418
rect 200620 283098 200652 283334
rect 200888 283098 200972 283334
rect 201208 283098 201240 283334
rect 236620 283418 236652 283654
rect 236888 283418 236972 283654
rect 237208 283418 237240 283654
rect 236620 283334 237240 283418
rect 236620 283098 236652 283334
rect 236888 283098 236972 283334
rect 237208 283098 237240 283334
rect 272620 283418 272652 283654
rect 272888 283418 272972 283654
rect 273208 283418 273240 283654
rect 272620 283334 273240 283418
rect 272620 283098 272652 283334
rect 272888 283098 272972 283334
rect 273208 283098 273240 283334
rect 308620 283418 308652 283654
rect 308888 283418 308972 283654
rect 309208 283418 309240 283654
rect 308620 283334 309240 283418
rect 308620 283098 308652 283334
rect 308888 283098 308972 283334
rect 309208 283098 309240 283334
rect 344620 283418 344652 283654
rect 344888 283418 344972 283654
rect 345208 283418 345240 283654
rect 344620 283334 345240 283418
rect 344620 283098 344652 283334
rect 344888 283098 344972 283334
rect 345208 283098 345240 283334
rect 380620 283418 380652 283654
rect 380888 283418 380972 283654
rect 381208 283418 381240 283654
rect 380620 283334 381240 283418
rect 380620 283098 380652 283334
rect 380888 283098 380972 283334
rect 381208 283098 381240 283334
rect 416620 283418 416652 283654
rect 416888 283418 416972 283654
rect 417208 283418 417240 283654
rect 416620 283334 417240 283418
rect 416620 283098 416652 283334
rect 416888 283098 416972 283334
rect 417208 283098 417240 283334
rect 452620 283418 452652 283654
rect 452888 283418 452972 283654
rect 453208 283418 453240 283654
rect 452620 283334 453240 283418
rect 452620 283098 452652 283334
rect 452888 283098 452972 283334
rect 453208 283098 453240 283334
rect 488620 283418 488652 283654
rect 488888 283418 488972 283654
rect 489208 283418 489240 283654
rect 488620 283334 489240 283418
rect 488620 283098 488652 283334
rect 488888 283098 488972 283334
rect 489208 283098 489240 283334
rect 524620 283418 524652 283654
rect 524888 283418 524972 283654
rect 525208 283418 525240 283654
rect 524620 283334 525240 283418
rect 524620 283098 524652 283334
rect 524888 283098 524972 283334
rect 525208 283098 525240 283334
rect 560620 283418 560652 283654
rect 560888 283418 560972 283654
rect 561208 283418 561240 283654
rect 560620 283334 561240 283418
rect 560620 283098 560652 283334
rect 560888 283098 560972 283334
rect 561208 283098 561240 283334
rect 570260 283418 570292 283654
rect 570528 283418 570612 283654
rect 570848 283418 570880 283654
rect 570260 283334 570880 283418
rect 570260 283098 570292 283334
rect 570528 283098 570612 283334
rect 570848 283098 570880 283334
rect -2006 243654 -1386 283098
rect 580594 262254 581214 301698
rect 580594 262018 580626 262254
rect 580862 262018 580946 262254
rect 581182 262018 581214 262254
rect 580594 261934 581214 262018
rect 580594 261698 580626 261934
rect 580862 261698 580946 261934
rect 581182 261698 581214 261934
rect 7844 247138 7876 247374
rect 8112 247138 8196 247374
rect 8432 247138 8464 247374
rect 7844 247054 8464 247138
rect 7844 246818 7876 247054
rect 8112 246818 8196 247054
rect 8432 246818 8464 247054
rect 38000 247138 38032 247374
rect 38268 247138 38352 247374
rect 38588 247138 38620 247374
rect 38000 247054 38620 247138
rect 38000 246818 38032 247054
rect 38268 246818 38352 247054
rect 38588 246818 38620 247054
rect 74000 247138 74032 247374
rect 74268 247138 74352 247374
rect 74588 247138 74620 247374
rect 74000 247054 74620 247138
rect 74000 246818 74032 247054
rect 74268 246818 74352 247054
rect 74588 246818 74620 247054
rect 110000 247138 110032 247374
rect 110268 247138 110352 247374
rect 110588 247138 110620 247374
rect 110000 247054 110620 247138
rect 110000 246818 110032 247054
rect 110268 246818 110352 247054
rect 110588 246818 110620 247054
rect 146000 247138 146032 247374
rect 146268 247138 146352 247374
rect 146588 247138 146620 247374
rect 146000 247054 146620 247138
rect 146000 246818 146032 247054
rect 146268 246818 146352 247054
rect 146588 246818 146620 247054
rect 182000 247138 182032 247374
rect 182268 247138 182352 247374
rect 182588 247138 182620 247374
rect 182000 247054 182620 247138
rect 182000 246818 182032 247054
rect 182268 246818 182352 247054
rect 182588 246818 182620 247054
rect 218000 247138 218032 247374
rect 218268 247138 218352 247374
rect 218588 247138 218620 247374
rect 218000 247054 218620 247138
rect 218000 246818 218032 247054
rect 218268 246818 218352 247054
rect 218588 246818 218620 247054
rect 254000 247138 254032 247374
rect 254268 247138 254352 247374
rect 254588 247138 254620 247374
rect 254000 247054 254620 247138
rect 254000 246818 254032 247054
rect 254268 246818 254352 247054
rect 254588 246818 254620 247054
rect 290000 247138 290032 247374
rect 290268 247138 290352 247374
rect 290588 247138 290620 247374
rect 290000 247054 290620 247138
rect 290000 246818 290032 247054
rect 290268 246818 290352 247054
rect 290588 246818 290620 247054
rect 326000 247138 326032 247374
rect 326268 247138 326352 247374
rect 326588 247138 326620 247374
rect 326000 247054 326620 247138
rect 326000 246818 326032 247054
rect 326268 246818 326352 247054
rect 326588 246818 326620 247054
rect 362000 247138 362032 247374
rect 362268 247138 362352 247374
rect 362588 247138 362620 247374
rect 362000 247054 362620 247138
rect 362000 246818 362032 247054
rect 362268 246818 362352 247054
rect 362588 246818 362620 247054
rect 398000 247138 398032 247374
rect 398268 247138 398352 247374
rect 398588 247138 398620 247374
rect 398000 247054 398620 247138
rect 398000 246818 398032 247054
rect 398268 246818 398352 247054
rect 398588 246818 398620 247054
rect 434000 247138 434032 247374
rect 434268 247138 434352 247374
rect 434588 247138 434620 247374
rect 434000 247054 434620 247138
rect 434000 246818 434032 247054
rect 434268 246818 434352 247054
rect 434588 246818 434620 247054
rect 470000 247138 470032 247374
rect 470268 247138 470352 247374
rect 470588 247138 470620 247374
rect 470000 247054 470620 247138
rect 470000 246818 470032 247054
rect 470268 246818 470352 247054
rect 470588 246818 470620 247054
rect 506000 247138 506032 247374
rect 506268 247138 506352 247374
rect 506588 247138 506620 247374
rect 506000 247054 506620 247138
rect 506000 246818 506032 247054
rect 506268 246818 506352 247054
rect 506588 246818 506620 247054
rect 542000 247138 542032 247374
rect 542268 247138 542352 247374
rect 542588 247138 542620 247374
rect 542000 247054 542620 247138
rect 542000 246818 542032 247054
rect 542268 246818 542352 247054
rect 542588 246818 542620 247054
rect 571500 247138 571532 247374
rect 571768 247138 571852 247374
rect 572088 247138 572120 247374
rect 571500 247054 572120 247138
rect 571500 246818 571532 247054
rect 571768 246818 571852 247054
rect 572088 246818 572120 247054
rect -2006 243418 -1974 243654
rect -1738 243418 -1654 243654
rect -1418 243418 -1386 243654
rect -2006 243334 -1386 243418
rect -2006 243098 -1974 243334
rect -1738 243098 -1654 243334
rect -1418 243098 -1386 243334
rect 9084 243418 9116 243654
rect 9352 243418 9436 243654
rect 9672 243418 9704 243654
rect 9084 243334 9704 243418
rect 9084 243098 9116 243334
rect 9352 243098 9436 243334
rect 9672 243098 9704 243334
rect 56620 243418 56652 243654
rect 56888 243418 56972 243654
rect 57208 243418 57240 243654
rect 56620 243334 57240 243418
rect 56620 243098 56652 243334
rect 56888 243098 56972 243334
rect 57208 243098 57240 243334
rect 92620 243418 92652 243654
rect 92888 243418 92972 243654
rect 93208 243418 93240 243654
rect 92620 243334 93240 243418
rect 92620 243098 92652 243334
rect 92888 243098 92972 243334
rect 93208 243098 93240 243334
rect 128620 243418 128652 243654
rect 128888 243418 128972 243654
rect 129208 243418 129240 243654
rect 128620 243334 129240 243418
rect 128620 243098 128652 243334
rect 128888 243098 128972 243334
rect 129208 243098 129240 243334
rect 164620 243418 164652 243654
rect 164888 243418 164972 243654
rect 165208 243418 165240 243654
rect 164620 243334 165240 243418
rect 164620 243098 164652 243334
rect 164888 243098 164972 243334
rect 165208 243098 165240 243334
rect 200620 243418 200652 243654
rect 200888 243418 200972 243654
rect 201208 243418 201240 243654
rect 200620 243334 201240 243418
rect 200620 243098 200652 243334
rect 200888 243098 200972 243334
rect 201208 243098 201240 243334
rect 236620 243418 236652 243654
rect 236888 243418 236972 243654
rect 237208 243418 237240 243654
rect 236620 243334 237240 243418
rect 236620 243098 236652 243334
rect 236888 243098 236972 243334
rect 237208 243098 237240 243334
rect 272620 243418 272652 243654
rect 272888 243418 272972 243654
rect 273208 243418 273240 243654
rect 272620 243334 273240 243418
rect 272620 243098 272652 243334
rect 272888 243098 272972 243334
rect 273208 243098 273240 243334
rect 308620 243418 308652 243654
rect 308888 243418 308972 243654
rect 309208 243418 309240 243654
rect 308620 243334 309240 243418
rect 308620 243098 308652 243334
rect 308888 243098 308972 243334
rect 309208 243098 309240 243334
rect 344620 243418 344652 243654
rect 344888 243418 344972 243654
rect 345208 243418 345240 243654
rect 344620 243334 345240 243418
rect 344620 243098 344652 243334
rect 344888 243098 344972 243334
rect 345208 243098 345240 243334
rect 380620 243418 380652 243654
rect 380888 243418 380972 243654
rect 381208 243418 381240 243654
rect 380620 243334 381240 243418
rect 380620 243098 380652 243334
rect 380888 243098 380972 243334
rect 381208 243098 381240 243334
rect 416620 243418 416652 243654
rect 416888 243418 416972 243654
rect 417208 243418 417240 243654
rect 416620 243334 417240 243418
rect 416620 243098 416652 243334
rect 416888 243098 416972 243334
rect 417208 243098 417240 243334
rect 452620 243418 452652 243654
rect 452888 243418 452972 243654
rect 453208 243418 453240 243654
rect 452620 243334 453240 243418
rect 452620 243098 452652 243334
rect 452888 243098 452972 243334
rect 453208 243098 453240 243334
rect 488620 243418 488652 243654
rect 488888 243418 488972 243654
rect 489208 243418 489240 243654
rect 488620 243334 489240 243418
rect 488620 243098 488652 243334
rect 488888 243098 488972 243334
rect 489208 243098 489240 243334
rect 524620 243418 524652 243654
rect 524888 243418 524972 243654
rect 525208 243418 525240 243654
rect 524620 243334 525240 243418
rect 524620 243098 524652 243334
rect 524888 243098 524972 243334
rect 525208 243098 525240 243334
rect 560620 243418 560652 243654
rect 560888 243418 560972 243654
rect 561208 243418 561240 243654
rect 560620 243334 561240 243418
rect 560620 243098 560652 243334
rect 560888 243098 560972 243334
rect 561208 243098 561240 243334
rect 570260 243418 570292 243654
rect 570528 243418 570612 243654
rect 570848 243418 570880 243654
rect 570260 243334 570880 243418
rect 570260 243098 570292 243334
rect 570528 243098 570612 243334
rect 570848 243098 570880 243334
rect -2006 203654 -1386 243098
rect 580594 222254 581214 261698
rect 580594 222018 580626 222254
rect 580862 222018 580946 222254
rect 581182 222018 581214 222254
rect 580594 221934 581214 222018
rect 580594 221698 580626 221934
rect 580862 221698 580946 221934
rect 581182 221698 581214 221934
rect 7844 207138 7876 207374
rect 8112 207138 8196 207374
rect 8432 207138 8464 207374
rect 7844 207054 8464 207138
rect 7844 206818 7876 207054
rect 8112 206818 8196 207054
rect 8432 206818 8464 207054
rect 38000 207138 38032 207374
rect 38268 207138 38352 207374
rect 38588 207138 38620 207374
rect 38000 207054 38620 207138
rect 38000 206818 38032 207054
rect 38268 206818 38352 207054
rect 38588 206818 38620 207054
rect 74000 207138 74032 207374
rect 74268 207138 74352 207374
rect 74588 207138 74620 207374
rect 74000 207054 74620 207138
rect 74000 206818 74032 207054
rect 74268 206818 74352 207054
rect 74588 206818 74620 207054
rect 110000 207138 110032 207374
rect 110268 207138 110352 207374
rect 110588 207138 110620 207374
rect 110000 207054 110620 207138
rect 110000 206818 110032 207054
rect 110268 206818 110352 207054
rect 110588 206818 110620 207054
rect 146000 207138 146032 207374
rect 146268 207138 146352 207374
rect 146588 207138 146620 207374
rect 146000 207054 146620 207138
rect 146000 206818 146032 207054
rect 146268 206818 146352 207054
rect 146588 206818 146620 207054
rect 182000 207138 182032 207374
rect 182268 207138 182352 207374
rect 182588 207138 182620 207374
rect 182000 207054 182620 207138
rect 182000 206818 182032 207054
rect 182268 206818 182352 207054
rect 182588 206818 182620 207054
rect 218000 207138 218032 207374
rect 218268 207138 218352 207374
rect 218588 207138 218620 207374
rect 218000 207054 218620 207138
rect 218000 206818 218032 207054
rect 218268 206818 218352 207054
rect 218588 206818 218620 207054
rect 254000 207138 254032 207374
rect 254268 207138 254352 207374
rect 254588 207138 254620 207374
rect 254000 207054 254620 207138
rect 254000 206818 254032 207054
rect 254268 206818 254352 207054
rect 254588 206818 254620 207054
rect 290000 207138 290032 207374
rect 290268 207138 290352 207374
rect 290588 207138 290620 207374
rect 290000 207054 290620 207138
rect 290000 206818 290032 207054
rect 290268 206818 290352 207054
rect 290588 206818 290620 207054
rect 326000 207138 326032 207374
rect 326268 207138 326352 207374
rect 326588 207138 326620 207374
rect 326000 207054 326620 207138
rect 326000 206818 326032 207054
rect 326268 206818 326352 207054
rect 326588 206818 326620 207054
rect 362000 207138 362032 207374
rect 362268 207138 362352 207374
rect 362588 207138 362620 207374
rect 362000 207054 362620 207138
rect 362000 206818 362032 207054
rect 362268 206818 362352 207054
rect 362588 206818 362620 207054
rect 398000 207138 398032 207374
rect 398268 207138 398352 207374
rect 398588 207138 398620 207374
rect 398000 207054 398620 207138
rect 398000 206818 398032 207054
rect 398268 206818 398352 207054
rect 398588 206818 398620 207054
rect 434000 207138 434032 207374
rect 434268 207138 434352 207374
rect 434588 207138 434620 207374
rect 434000 207054 434620 207138
rect 434000 206818 434032 207054
rect 434268 206818 434352 207054
rect 434588 206818 434620 207054
rect 470000 207138 470032 207374
rect 470268 207138 470352 207374
rect 470588 207138 470620 207374
rect 470000 207054 470620 207138
rect 470000 206818 470032 207054
rect 470268 206818 470352 207054
rect 470588 206818 470620 207054
rect 506000 207138 506032 207374
rect 506268 207138 506352 207374
rect 506588 207138 506620 207374
rect 506000 207054 506620 207138
rect 506000 206818 506032 207054
rect 506268 206818 506352 207054
rect 506588 206818 506620 207054
rect 542000 207138 542032 207374
rect 542268 207138 542352 207374
rect 542588 207138 542620 207374
rect 542000 207054 542620 207138
rect 542000 206818 542032 207054
rect 542268 206818 542352 207054
rect 542588 206818 542620 207054
rect 571500 207138 571532 207374
rect 571768 207138 571852 207374
rect 572088 207138 572120 207374
rect 571500 207054 572120 207138
rect 571500 206818 571532 207054
rect 571768 206818 571852 207054
rect 572088 206818 572120 207054
rect -2006 203418 -1974 203654
rect -1738 203418 -1654 203654
rect -1418 203418 -1386 203654
rect -2006 203334 -1386 203418
rect -2006 203098 -1974 203334
rect -1738 203098 -1654 203334
rect -1418 203098 -1386 203334
rect 9084 203418 9116 203654
rect 9352 203418 9436 203654
rect 9672 203418 9704 203654
rect 9084 203334 9704 203418
rect 9084 203098 9116 203334
rect 9352 203098 9436 203334
rect 9672 203098 9704 203334
rect 56620 203418 56652 203654
rect 56888 203418 56972 203654
rect 57208 203418 57240 203654
rect 56620 203334 57240 203418
rect 56620 203098 56652 203334
rect 56888 203098 56972 203334
rect 57208 203098 57240 203334
rect 92620 203418 92652 203654
rect 92888 203418 92972 203654
rect 93208 203418 93240 203654
rect 92620 203334 93240 203418
rect 92620 203098 92652 203334
rect 92888 203098 92972 203334
rect 93208 203098 93240 203334
rect 128620 203418 128652 203654
rect 128888 203418 128972 203654
rect 129208 203418 129240 203654
rect 128620 203334 129240 203418
rect 128620 203098 128652 203334
rect 128888 203098 128972 203334
rect 129208 203098 129240 203334
rect 164620 203418 164652 203654
rect 164888 203418 164972 203654
rect 165208 203418 165240 203654
rect 164620 203334 165240 203418
rect 164620 203098 164652 203334
rect 164888 203098 164972 203334
rect 165208 203098 165240 203334
rect 200620 203418 200652 203654
rect 200888 203418 200972 203654
rect 201208 203418 201240 203654
rect 200620 203334 201240 203418
rect 200620 203098 200652 203334
rect 200888 203098 200972 203334
rect 201208 203098 201240 203334
rect 236620 203418 236652 203654
rect 236888 203418 236972 203654
rect 237208 203418 237240 203654
rect 236620 203334 237240 203418
rect 236620 203098 236652 203334
rect 236888 203098 236972 203334
rect 237208 203098 237240 203334
rect 272620 203418 272652 203654
rect 272888 203418 272972 203654
rect 273208 203418 273240 203654
rect 272620 203334 273240 203418
rect 272620 203098 272652 203334
rect 272888 203098 272972 203334
rect 273208 203098 273240 203334
rect 308620 203418 308652 203654
rect 308888 203418 308972 203654
rect 309208 203418 309240 203654
rect 308620 203334 309240 203418
rect 308620 203098 308652 203334
rect 308888 203098 308972 203334
rect 309208 203098 309240 203334
rect 344620 203418 344652 203654
rect 344888 203418 344972 203654
rect 345208 203418 345240 203654
rect 344620 203334 345240 203418
rect 344620 203098 344652 203334
rect 344888 203098 344972 203334
rect 345208 203098 345240 203334
rect 380620 203418 380652 203654
rect 380888 203418 380972 203654
rect 381208 203418 381240 203654
rect 380620 203334 381240 203418
rect 380620 203098 380652 203334
rect 380888 203098 380972 203334
rect 381208 203098 381240 203334
rect 416620 203418 416652 203654
rect 416888 203418 416972 203654
rect 417208 203418 417240 203654
rect 416620 203334 417240 203418
rect 416620 203098 416652 203334
rect 416888 203098 416972 203334
rect 417208 203098 417240 203334
rect 452620 203418 452652 203654
rect 452888 203418 452972 203654
rect 453208 203418 453240 203654
rect 452620 203334 453240 203418
rect 452620 203098 452652 203334
rect 452888 203098 452972 203334
rect 453208 203098 453240 203334
rect 488620 203418 488652 203654
rect 488888 203418 488972 203654
rect 489208 203418 489240 203654
rect 488620 203334 489240 203418
rect 488620 203098 488652 203334
rect 488888 203098 488972 203334
rect 489208 203098 489240 203334
rect 524620 203418 524652 203654
rect 524888 203418 524972 203654
rect 525208 203418 525240 203654
rect 524620 203334 525240 203418
rect 524620 203098 524652 203334
rect 524888 203098 524972 203334
rect 525208 203098 525240 203334
rect 560620 203418 560652 203654
rect 560888 203418 560972 203654
rect 561208 203418 561240 203654
rect 560620 203334 561240 203418
rect 560620 203098 560652 203334
rect 560888 203098 560972 203334
rect 561208 203098 561240 203334
rect 570260 203418 570292 203654
rect 570528 203418 570612 203654
rect 570848 203418 570880 203654
rect 570260 203334 570880 203418
rect 570260 203098 570292 203334
rect 570528 203098 570612 203334
rect 570848 203098 570880 203334
rect -2006 163654 -1386 203098
rect 580594 182254 581214 221698
rect 580594 182018 580626 182254
rect 580862 182018 580946 182254
rect 581182 182018 581214 182254
rect 580594 181934 581214 182018
rect 580594 181698 580626 181934
rect 580862 181698 580946 181934
rect 581182 181698 581214 181934
rect 60560 167374 60920 167406
rect 7844 167138 7876 167374
rect 8112 167138 8196 167374
rect 8432 167138 8464 167374
rect 7844 167054 8464 167138
rect 7844 166818 7876 167054
rect 8112 166818 8196 167054
rect 8432 166818 8464 167054
rect 38000 167138 38032 167374
rect 38268 167138 38352 167374
rect 38588 167138 38620 167374
rect 38000 167054 38620 167138
rect 38000 166818 38032 167054
rect 38268 166818 38352 167054
rect 38588 166818 38620 167054
rect 60560 167138 60622 167374
rect 60858 167138 60920 167374
rect 60560 167054 60920 167138
rect 60560 166818 60622 167054
rect 60858 166818 60920 167054
rect 60560 166786 60920 166818
rect 159036 167374 159396 167406
rect 185560 167374 185920 167406
rect 159036 167138 159098 167374
rect 159334 167138 159396 167374
rect 159036 167054 159396 167138
rect 159036 166818 159098 167054
rect 159334 166818 159396 167054
rect 182000 167138 182032 167374
rect 182268 167138 182352 167374
rect 182588 167138 182620 167374
rect 182000 167054 182620 167138
rect 182000 166818 182032 167054
rect 182268 166818 182352 167054
rect 182588 166818 182620 167054
rect 185560 167138 185622 167374
rect 185858 167138 185920 167374
rect 185560 167054 185920 167138
rect 185560 166818 185622 167054
rect 185858 166818 185920 167054
rect 159036 166786 159396 166818
rect 185560 166786 185920 166818
rect 284036 167374 284396 167406
rect 310560 167374 310920 167406
rect 284036 167138 284098 167374
rect 284334 167138 284396 167374
rect 284036 167054 284396 167138
rect 284036 166818 284098 167054
rect 284334 166818 284396 167054
rect 290000 167138 290032 167374
rect 290268 167138 290352 167374
rect 290588 167138 290620 167374
rect 290000 167054 290620 167138
rect 290000 166818 290032 167054
rect 290268 166818 290352 167054
rect 290588 166818 290620 167054
rect 310560 167138 310622 167374
rect 310858 167138 310920 167374
rect 310560 167054 310920 167138
rect 310560 166818 310622 167054
rect 310858 166818 310920 167054
rect 284036 166786 284396 166818
rect 310560 166786 310920 166818
rect 409036 167374 409396 167406
rect 436560 167374 436920 167406
rect 409036 167138 409098 167374
rect 409334 167138 409396 167374
rect 409036 167054 409396 167138
rect 409036 166818 409098 167054
rect 409334 166818 409396 167054
rect 434000 167138 434032 167374
rect 434268 167138 434352 167374
rect 434588 167138 434620 167374
rect 434000 167054 434620 167138
rect 434000 166818 434032 167054
rect 434268 166818 434352 167054
rect 434588 166818 434620 167054
rect 436560 167138 436622 167374
rect 436858 167138 436920 167374
rect 436560 167054 436920 167138
rect 436560 166818 436622 167054
rect 436858 166818 436920 167054
rect 409036 166786 409396 166818
rect 436560 166786 436920 166818
rect 535036 167374 535396 167406
rect 535036 167138 535098 167374
rect 535334 167138 535396 167374
rect 535036 167054 535396 167138
rect 535036 166818 535098 167054
rect 535334 166818 535396 167054
rect 542000 167138 542032 167374
rect 542268 167138 542352 167374
rect 542588 167138 542620 167374
rect 542000 167054 542620 167138
rect 542000 166818 542032 167054
rect 542268 166818 542352 167054
rect 542588 166818 542620 167054
rect 571500 167138 571532 167374
rect 571768 167138 571852 167374
rect 572088 167138 572120 167374
rect 571500 167054 572120 167138
rect 571500 166818 571532 167054
rect 571768 166818 571852 167054
rect 572088 166818 572120 167054
rect 535036 166786 535396 166818
rect 61280 163654 61640 163686
rect -2006 163418 -1974 163654
rect -1738 163418 -1654 163654
rect -1418 163418 -1386 163654
rect -2006 163334 -1386 163418
rect -2006 163098 -1974 163334
rect -1738 163098 -1654 163334
rect -1418 163098 -1386 163334
rect 9084 163418 9116 163654
rect 9352 163418 9436 163654
rect 9672 163418 9704 163654
rect 9084 163334 9704 163418
rect 9084 163098 9116 163334
rect 9352 163098 9436 163334
rect 9672 163098 9704 163334
rect 56620 163418 56652 163654
rect 56888 163418 56972 163654
rect 57208 163418 57240 163654
rect 56620 163334 57240 163418
rect 56620 163098 56652 163334
rect 56888 163098 56972 163334
rect 57208 163098 57240 163334
rect 61280 163418 61342 163654
rect 61578 163418 61640 163654
rect 61280 163334 61640 163418
rect 61280 163098 61342 163334
rect 61578 163098 61640 163334
rect -2006 123654 -1386 163098
rect 61280 163066 61640 163098
rect 158316 163654 158676 163686
rect 186280 163654 186640 163686
rect 158316 163418 158378 163654
rect 158614 163418 158676 163654
rect 158316 163334 158676 163418
rect 158316 163098 158378 163334
rect 158614 163098 158676 163334
rect 164620 163418 164652 163654
rect 164888 163418 164972 163654
rect 165208 163418 165240 163654
rect 164620 163334 165240 163418
rect 164620 163098 164652 163334
rect 164888 163098 164972 163334
rect 165208 163098 165240 163334
rect 186280 163418 186342 163654
rect 186578 163418 186640 163654
rect 186280 163334 186640 163418
rect 186280 163098 186342 163334
rect 186578 163098 186640 163334
rect 158316 163066 158676 163098
rect 186280 163066 186640 163098
rect 283316 163654 283676 163686
rect 311280 163654 311640 163686
rect 283316 163418 283378 163654
rect 283614 163418 283676 163654
rect 283316 163334 283676 163418
rect 283316 163098 283378 163334
rect 283614 163098 283676 163334
rect 308620 163418 308652 163654
rect 308888 163418 308972 163654
rect 309208 163418 309240 163654
rect 308620 163334 309240 163418
rect 308620 163098 308652 163334
rect 308888 163098 308972 163334
rect 309208 163098 309240 163334
rect 311280 163418 311342 163654
rect 311578 163418 311640 163654
rect 311280 163334 311640 163418
rect 311280 163098 311342 163334
rect 311578 163098 311640 163334
rect 283316 163066 283676 163098
rect 311280 163066 311640 163098
rect 408316 163654 408676 163686
rect 437280 163654 437640 163686
rect 408316 163418 408378 163654
rect 408614 163418 408676 163654
rect 408316 163334 408676 163418
rect 408316 163098 408378 163334
rect 408614 163098 408676 163334
rect 416620 163418 416652 163654
rect 416888 163418 416972 163654
rect 417208 163418 417240 163654
rect 416620 163334 417240 163418
rect 416620 163098 416652 163334
rect 416888 163098 416972 163334
rect 417208 163098 417240 163334
rect 437280 163418 437342 163654
rect 437578 163418 437640 163654
rect 437280 163334 437640 163418
rect 437280 163098 437342 163334
rect 437578 163098 437640 163334
rect 408316 163066 408676 163098
rect 437280 163066 437640 163098
rect 534316 163654 534676 163686
rect 534316 163418 534378 163654
rect 534614 163418 534676 163654
rect 534316 163334 534676 163418
rect 534316 163098 534378 163334
rect 534614 163098 534676 163334
rect 560620 163418 560652 163654
rect 560888 163418 560972 163654
rect 561208 163418 561240 163654
rect 560620 163334 561240 163418
rect 560620 163098 560652 163334
rect 560888 163098 560972 163334
rect 561208 163098 561240 163334
rect 570260 163418 570292 163654
rect 570528 163418 570612 163654
rect 570848 163418 570880 163654
rect 570260 163334 570880 163418
rect 570260 163098 570292 163334
rect 570528 163098 570612 163334
rect 570848 163098 570880 163334
rect 534316 163066 534676 163098
rect 580594 142254 581214 181698
rect 580594 142018 580626 142254
rect 580862 142018 580946 142254
rect 581182 142018 581214 142254
rect 580594 141934 581214 142018
rect 580594 141698 580626 141934
rect 580862 141698 580946 141934
rect 581182 141698 581214 141934
rect 60560 127374 60920 127406
rect 7844 127138 7876 127374
rect 8112 127138 8196 127374
rect 8432 127138 8464 127374
rect 7844 127054 8464 127138
rect 7844 126818 7876 127054
rect 8112 126818 8196 127054
rect 8432 126818 8464 127054
rect 38000 127138 38032 127374
rect 38268 127138 38352 127374
rect 38588 127138 38620 127374
rect 38000 127054 38620 127138
rect 38000 126818 38032 127054
rect 38268 126818 38352 127054
rect 38588 126818 38620 127054
rect 60560 127138 60622 127374
rect 60858 127138 60920 127374
rect 60560 127054 60920 127138
rect 60560 126818 60622 127054
rect 60858 126818 60920 127054
rect 60560 126786 60920 126818
rect 159036 127374 159396 127406
rect 185560 127374 185920 127406
rect 159036 127138 159098 127374
rect 159334 127138 159396 127374
rect 159036 127054 159396 127138
rect 159036 126818 159098 127054
rect 159334 126818 159396 127054
rect 182000 127138 182032 127374
rect 182268 127138 182352 127374
rect 182588 127138 182620 127374
rect 182000 127054 182620 127138
rect 182000 126818 182032 127054
rect 182268 126818 182352 127054
rect 182588 126818 182620 127054
rect 185560 127138 185622 127374
rect 185858 127138 185920 127374
rect 185560 127054 185920 127138
rect 185560 126818 185622 127054
rect 185858 126818 185920 127054
rect 159036 126786 159396 126818
rect 185560 126786 185920 126818
rect 284036 127374 284396 127406
rect 310560 127374 310920 127406
rect 284036 127138 284098 127374
rect 284334 127138 284396 127374
rect 284036 127054 284396 127138
rect 284036 126818 284098 127054
rect 284334 126818 284396 127054
rect 290000 127138 290032 127374
rect 290268 127138 290352 127374
rect 290588 127138 290620 127374
rect 290000 127054 290620 127138
rect 290000 126818 290032 127054
rect 290268 126818 290352 127054
rect 290588 126818 290620 127054
rect 310560 127138 310622 127374
rect 310858 127138 310920 127374
rect 310560 127054 310920 127138
rect 310560 126818 310622 127054
rect 310858 126818 310920 127054
rect 284036 126786 284396 126818
rect 310560 126786 310920 126818
rect 409036 127374 409396 127406
rect 436560 127374 436920 127406
rect 409036 127138 409098 127374
rect 409334 127138 409396 127374
rect 409036 127054 409396 127138
rect 409036 126818 409098 127054
rect 409334 126818 409396 127054
rect 434000 127138 434032 127374
rect 434268 127138 434352 127374
rect 434588 127138 434620 127374
rect 434000 127054 434620 127138
rect 434000 126818 434032 127054
rect 434268 126818 434352 127054
rect 434588 126818 434620 127054
rect 436560 127138 436622 127374
rect 436858 127138 436920 127374
rect 436560 127054 436920 127138
rect 436560 126818 436622 127054
rect 436858 126818 436920 127054
rect 409036 126786 409396 126818
rect 436560 126786 436920 126818
rect 535036 127374 535396 127406
rect 535036 127138 535098 127374
rect 535334 127138 535396 127374
rect 535036 127054 535396 127138
rect 535036 126818 535098 127054
rect 535334 126818 535396 127054
rect 542000 127138 542032 127374
rect 542268 127138 542352 127374
rect 542588 127138 542620 127374
rect 542000 127054 542620 127138
rect 542000 126818 542032 127054
rect 542268 126818 542352 127054
rect 542588 126818 542620 127054
rect 571500 127138 571532 127374
rect 571768 127138 571852 127374
rect 572088 127138 572120 127374
rect 571500 127054 572120 127138
rect 571500 126818 571532 127054
rect 571768 126818 571852 127054
rect 572088 126818 572120 127054
rect 535036 126786 535396 126818
rect 61280 123654 61640 123686
rect -2006 123418 -1974 123654
rect -1738 123418 -1654 123654
rect -1418 123418 -1386 123654
rect -2006 123334 -1386 123418
rect -2006 123098 -1974 123334
rect -1738 123098 -1654 123334
rect -1418 123098 -1386 123334
rect 9084 123418 9116 123654
rect 9352 123418 9436 123654
rect 9672 123418 9704 123654
rect 9084 123334 9704 123418
rect 9084 123098 9116 123334
rect 9352 123098 9436 123334
rect 9672 123098 9704 123334
rect 56620 123418 56652 123654
rect 56888 123418 56972 123654
rect 57208 123418 57240 123654
rect 56620 123334 57240 123418
rect 56620 123098 56652 123334
rect 56888 123098 56972 123334
rect 57208 123098 57240 123334
rect 61280 123418 61342 123654
rect 61578 123418 61640 123654
rect 61280 123334 61640 123418
rect 61280 123098 61342 123334
rect 61578 123098 61640 123334
rect -2006 83654 -1386 123098
rect 61280 123066 61640 123098
rect 158316 123654 158676 123686
rect 186280 123654 186640 123686
rect 158316 123418 158378 123654
rect 158614 123418 158676 123654
rect 158316 123334 158676 123418
rect 158316 123098 158378 123334
rect 158614 123098 158676 123334
rect 164620 123418 164652 123654
rect 164888 123418 164972 123654
rect 165208 123418 165240 123654
rect 164620 123334 165240 123418
rect 164620 123098 164652 123334
rect 164888 123098 164972 123334
rect 165208 123098 165240 123334
rect 186280 123418 186342 123654
rect 186578 123418 186640 123654
rect 186280 123334 186640 123418
rect 186280 123098 186342 123334
rect 186578 123098 186640 123334
rect 158316 123066 158676 123098
rect 186280 123066 186640 123098
rect 283316 123654 283676 123686
rect 311280 123654 311640 123686
rect 283316 123418 283378 123654
rect 283614 123418 283676 123654
rect 283316 123334 283676 123418
rect 283316 123098 283378 123334
rect 283614 123098 283676 123334
rect 308620 123418 308652 123654
rect 308888 123418 308972 123654
rect 309208 123418 309240 123654
rect 308620 123334 309240 123418
rect 308620 123098 308652 123334
rect 308888 123098 308972 123334
rect 309208 123098 309240 123334
rect 311280 123418 311342 123654
rect 311578 123418 311640 123654
rect 311280 123334 311640 123418
rect 311280 123098 311342 123334
rect 311578 123098 311640 123334
rect 283316 123066 283676 123098
rect 311280 123066 311640 123098
rect 408316 123654 408676 123686
rect 437280 123654 437640 123686
rect 408316 123418 408378 123654
rect 408614 123418 408676 123654
rect 408316 123334 408676 123418
rect 408316 123098 408378 123334
rect 408614 123098 408676 123334
rect 416620 123418 416652 123654
rect 416888 123418 416972 123654
rect 417208 123418 417240 123654
rect 416620 123334 417240 123418
rect 416620 123098 416652 123334
rect 416888 123098 416972 123334
rect 417208 123098 417240 123334
rect 437280 123418 437342 123654
rect 437578 123418 437640 123654
rect 437280 123334 437640 123418
rect 437280 123098 437342 123334
rect 437578 123098 437640 123334
rect 408316 123066 408676 123098
rect 437280 123066 437640 123098
rect 534316 123654 534676 123686
rect 534316 123418 534378 123654
rect 534614 123418 534676 123654
rect 534316 123334 534676 123418
rect 534316 123098 534378 123334
rect 534614 123098 534676 123334
rect 560620 123418 560652 123654
rect 560888 123418 560972 123654
rect 561208 123418 561240 123654
rect 560620 123334 561240 123418
rect 560620 123098 560652 123334
rect 560888 123098 560972 123334
rect 561208 123098 561240 123334
rect 570260 123418 570292 123654
rect 570528 123418 570612 123654
rect 570848 123418 570880 123654
rect 570260 123334 570880 123418
rect 570260 123098 570292 123334
rect 570528 123098 570612 123334
rect 570848 123098 570880 123334
rect 534316 123066 534676 123098
rect 61280 121244 61640 121300
rect 61280 121008 61342 121244
rect 61578 121008 61640 121244
rect 61280 120952 61640 121008
rect 62952 121244 63300 121300
rect 62952 121008 63008 121244
rect 63244 121008 63300 121244
rect 62952 120952 63300 121008
rect 281656 121244 282004 121300
rect 281656 121008 281712 121244
rect 281948 121008 282004 121244
rect 281656 120952 282004 121008
rect 283316 121244 283676 121300
rect 283316 121008 283378 121244
rect 283614 121008 283676 121244
rect 283316 120952 283676 121008
rect 311280 121244 311640 121300
rect 311280 121008 311342 121244
rect 311578 121008 311640 121244
rect 311280 120952 311640 121008
rect 312952 121244 313300 121300
rect 312952 121008 313008 121244
rect 313244 121008 313300 121244
rect 312952 120952 313300 121008
rect 532656 121244 533004 121300
rect 532656 121008 532712 121244
rect 532948 121008 533004 121244
rect 532656 120952 533004 121008
rect 534316 121244 534676 121300
rect 534316 121008 534378 121244
rect 534614 121008 534676 121244
rect 534316 120952 534676 121008
rect 157336 120564 157684 120620
rect 157336 120328 157392 120564
rect 157628 120328 157684 120564
rect 157336 120272 157684 120328
rect 159036 120564 159396 120620
rect 159036 120328 159098 120564
rect 159334 120328 159396 120564
rect 159036 120272 159396 120328
rect 185560 120564 185920 120620
rect 185560 120328 185622 120564
rect 185858 120328 185920 120564
rect 185560 120272 185920 120328
rect 187272 120564 187620 120620
rect 187272 120328 187328 120564
rect 187564 120328 187620 120564
rect 187272 120272 187620 120328
rect 407336 120564 407684 120620
rect 407336 120328 407392 120564
rect 407628 120328 407684 120564
rect 407336 120272 407684 120328
rect 409036 120564 409396 120620
rect 409036 120328 409098 120564
rect 409334 120328 409396 120564
rect 409036 120272 409396 120328
rect 436560 120564 436920 120620
rect 436560 120328 436622 120564
rect 436858 120328 436920 120564
rect 436560 120272 436920 120328
rect 438272 120564 438620 120620
rect 438272 120328 438328 120564
rect 438564 120328 438620 120564
rect 438272 120272 438620 120328
rect 580594 102254 581214 141698
rect 580594 102018 580626 102254
rect 580862 102018 580946 102254
rect 581182 102018 581214 102254
rect 580594 101934 581214 102018
rect 580594 101698 580626 101934
rect 580862 101698 580946 101934
rect 581182 101698 581214 101934
rect 60560 87374 60920 87406
rect 7844 87138 7876 87374
rect 8112 87138 8196 87374
rect 8432 87138 8464 87374
rect 7844 87054 8464 87138
rect 7844 86818 7876 87054
rect 8112 86818 8196 87054
rect 8432 86818 8464 87054
rect 38000 87138 38032 87374
rect 38268 87138 38352 87374
rect 38588 87138 38620 87374
rect 38000 87054 38620 87138
rect 38000 86818 38032 87054
rect 38268 86818 38352 87054
rect 38588 86818 38620 87054
rect 60560 87138 60622 87374
rect 60858 87138 60920 87374
rect 60560 87054 60920 87138
rect 60560 86818 60622 87054
rect 60858 86818 60920 87054
rect 60560 86786 60920 86818
rect 159036 87374 159396 87406
rect 185560 87374 185920 87406
rect 159036 87138 159098 87374
rect 159334 87138 159396 87374
rect 159036 87054 159396 87138
rect 159036 86818 159098 87054
rect 159334 86818 159396 87054
rect 182000 87138 182032 87374
rect 182268 87138 182352 87374
rect 182588 87138 182620 87374
rect 182000 87054 182620 87138
rect 182000 86818 182032 87054
rect 182268 86818 182352 87054
rect 182588 86818 182620 87054
rect 185560 87138 185622 87374
rect 185858 87138 185920 87374
rect 185560 87054 185920 87138
rect 185560 86818 185622 87054
rect 185858 86818 185920 87054
rect 159036 86786 159396 86818
rect 185560 86786 185920 86818
rect 284036 87374 284396 87406
rect 310560 87374 310920 87406
rect 284036 87138 284098 87374
rect 284334 87138 284396 87374
rect 284036 87054 284396 87138
rect 284036 86818 284098 87054
rect 284334 86818 284396 87054
rect 290000 87138 290032 87374
rect 290268 87138 290352 87374
rect 290588 87138 290620 87374
rect 290000 87054 290620 87138
rect 290000 86818 290032 87054
rect 290268 86818 290352 87054
rect 290588 86818 290620 87054
rect 310560 87138 310622 87374
rect 310858 87138 310920 87374
rect 310560 87054 310920 87138
rect 310560 86818 310622 87054
rect 310858 86818 310920 87054
rect 284036 86786 284396 86818
rect 310560 86786 310920 86818
rect 409036 87374 409396 87406
rect 436560 87374 436920 87406
rect 409036 87138 409098 87374
rect 409334 87138 409396 87374
rect 409036 87054 409396 87138
rect 409036 86818 409098 87054
rect 409334 86818 409396 87054
rect 434000 87138 434032 87374
rect 434268 87138 434352 87374
rect 434588 87138 434620 87374
rect 434000 87054 434620 87138
rect 434000 86818 434032 87054
rect 434268 86818 434352 87054
rect 434588 86818 434620 87054
rect 436560 87138 436622 87374
rect 436858 87138 436920 87374
rect 436560 87054 436920 87138
rect 436560 86818 436622 87054
rect 436858 86818 436920 87054
rect 409036 86786 409396 86818
rect 436560 86786 436920 86818
rect 535036 87374 535396 87406
rect 535036 87138 535098 87374
rect 535334 87138 535396 87374
rect 535036 87054 535396 87138
rect 535036 86818 535098 87054
rect 535334 86818 535396 87054
rect 542000 87138 542032 87374
rect 542268 87138 542352 87374
rect 542588 87138 542620 87374
rect 542000 87054 542620 87138
rect 542000 86818 542032 87054
rect 542268 86818 542352 87054
rect 542588 86818 542620 87054
rect 571500 87138 571532 87374
rect 571768 87138 571852 87374
rect 572088 87138 572120 87374
rect 571500 87054 572120 87138
rect 571500 86818 571532 87054
rect 571768 86818 571852 87054
rect 572088 86818 572120 87054
rect 535036 86786 535396 86818
rect 61280 83654 61640 83686
rect -2006 83418 -1974 83654
rect -1738 83418 -1654 83654
rect -1418 83418 -1386 83654
rect -2006 83334 -1386 83418
rect -2006 83098 -1974 83334
rect -1738 83098 -1654 83334
rect -1418 83098 -1386 83334
rect 9084 83418 9116 83654
rect 9352 83418 9436 83654
rect 9672 83418 9704 83654
rect 9084 83334 9704 83418
rect 9084 83098 9116 83334
rect 9352 83098 9436 83334
rect 9672 83098 9704 83334
rect 56620 83418 56652 83654
rect 56888 83418 56972 83654
rect 57208 83418 57240 83654
rect 56620 83334 57240 83418
rect 56620 83098 56652 83334
rect 56888 83098 56972 83334
rect 57208 83098 57240 83334
rect 61280 83418 61342 83654
rect 61578 83418 61640 83654
rect 61280 83334 61640 83418
rect 61280 83098 61342 83334
rect 61578 83098 61640 83334
rect -2006 43654 -1386 83098
rect 61280 83066 61640 83098
rect 158316 83654 158676 83686
rect 186280 83654 186640 83686
rect 158316 83418 158378 83654
rect 158614 83418 158676 83654
rect 158316 83334 158676 83418
rect 158316 83098 158378 83334
rect 158614 83098 158676 83334
rect 164620 83418 164652 83654
rect 164888 83418 164972 83654
rect 165208 83418 165240 83654
rect 164620 83334 165240 83418
rect 164620 83098 164652 83334
rect 164888 83098 164972 83334
rect 165208 83098 165240 83334
rect 186280 83418 186342 83654
rect 186578 83418 186640 83654
rect 186280 83334 186640 83418
rect 186280 83098 186342 83334
rect 186578 83098 186640 83334
rect 158316 83066 158676 83098
rect 186280 83066 186640 83098
rect 283316 83654 283676 83686
rect 311280 83654 311640 83686
rect 283316 83418 283378 83654
rect 283614 83418 283676 83654
rect 283316 83334 283676 83418
rect 283316 83098 283378 83334
rect 283614 83098 283676 83334
rect 308620 83418 308652 83654
rect 308888 83418 308972 83654
rect 309208 83418 309240 83654
rect 308620 83334 309240 83418
rect 308620 83098 308652 83334
rect 308888 83098 308972 83334
rect 309208 83098 309240 83334
rect 311280 83418 311342 83654
rect 311578 83418 311640 83654
rect 311280 83334 311640 83418
rect 311280 83098 311342 83334
rect 311578 83098 311640 83334
rect 283316 83066 283676 83098
rect 311280 83066 311640 83098
rect 408316 83654 408676 83686
rect 437280 83654 437640 83686
rect 408316 83418 408378 83654
rect 408614 83418 408676 83654
rect 408316 83334 408676 83418
rect 408316 83098 408378 83334
rect 408614 83098 408676 83334
rect 416620 83418 416652 83654
rect 416888 83418 416972 83654
rect 417208 83418 417240 83654
rect 416620 83334 417240 83418
rect 416620 83098 416652 83334
rect 416888 83098 416972 83334
rect 417208 83098 417240 83334
rect 437280 83418 437342 83654
rect 437578 83418 437640 83654
rect 437280 83334 437640 83418
rect 437280 83098 437342 83334
rect 437578 83098 437640 83334
rect 408316 83066 408676 83098
rect 437280 83066 437640 83098
rect 534316 83654 534676 83686
rect 534316 83418 534378 83654
rect 534614 83418 534676 83654
rect 534316 83334 534676 83418
rect 534316 83098 534378 83334
rect 534614 83098 534676 83334
rect 560620 83418 560652 83654
rect 560888 83418 560972 83654
rect 561208 83418 561240 83654
rect 560620 83334 561240 83418
rect 560620 83098 560652 83334
rect 560888 83098 560972 83334
rect 561208 83098 561240 83334
rect 570260 83418 570292 83654
rect 570528 83418 570612 83654
rect 570848 83418 570880 83654
rect 570260 83334 570880 83418
rect 570260 83098 570292 83334
rect 570528 83098 570612 83334
rect 570848 83098 570880 83334
rect 534316 83066 534676 83098
rect 580594 62254 581214 101698
rect 580594 62018 580626 62254
rect 580862 62018 580946 62254
rect 581182 62018 581214 62254
rect 580594 61934 581214 62018
rect 580594 61698 580626 61934
rect 580862 61698 580946 61934
rect 581182 61698 581214 61934
rect 60560 47374 60920 47406
rect 7844 47138 7876 47374
rect 8112 47138 8196 47374
rect 8432 47138 8464 47374
rect 7844 47054 8464 47138
rect 7844 46818 7876 47054
rect 8112 46818 8196 47054
rect 8432 46818 8464 47054
rect 38000 47138 38032 47374
rect 38268 47138 38352 47374
rect 38588 47138 38620 47374
rect 38000 47054 38620 47138
rect 38000 46818 38032 47054
rect 38268 46818 38352 47054
rect 38588 46818 38620 47054
rect 60560 47138 60622 47374
rect 60858 47138 60920 47374
rect 60560 47054 60920 47138
rect 60560 46818 60622 47054
rect 60858 46818 60920 47054
rect 60560 46786 60920 46818
rect 159036 47374 159396 47406
rect 185560 47374 185920 47406
rect 159036 47138 159098 47374
rect 159334 47138 159396 47374
rect 159036 47054 159396 47138
rect 159036 46818 159098 47054
rect 159334 46818 159396 47054
rect 182000 47138 182032 47374
rect 182268 47138 182352 47374
rect 182588 47138 182620 47374
rect 182000 47054 182620 47138
rect 182000 46818 182032 47054
rect 182268 46818 182352 47054
rect 182588 46818 182620 47054
rect 185560 47138 185622 47374
rect 185858 47138 185920 47374
rect 185560 47054 185920 47138
rect 185560 46818 185622 47054
rect 185858 46818 185920 47054
rect 159036 46786 159396 46818
rect 185560 46786 185920 46818
rect 284036 47374 284396 47406
rect 310560 47374 310920 47406
rect 284036 47138 284098 47374
rect 284334 47138 284396 47374
rect 284036 47054 284396 47138
rect 284036 46818 284098 47054
rect 284334 46818 284396 47054
rect 290000 47138 290032 47374
rect 290268 47138 290352 47374
rect 290588 47138 290620 47374
rect 290000 47054 290620 47138
rect 290000 46818 290032 47054
rect 290268 46818 290352 47054
rect 290588 46818 290620 47054
rect 310560 47138 310622 47374
rect 310858 47138 310920 47374
rect 310560 47054 310920 47138
rect 310560 46818 310622 47054
rect 310858 46818 310920 47054
rect 284036 46786 284396 46818
rect 310560 46786 310920 46818
rect 409036 47374 409396 47406
rect 436560 47374 436920 47406
rect 409036 47138 409098 47374
rect 409334 47138 409396 47374
rect 409036 47054 409396 47138
rect 409036 46818 409098 47054
rect 409334 46818 409396 47054
rect 434000 47138 434032 47374
rect 434268 47138 434352 47374
rect 434588 47138 434620 47374
rect 434000 47054 434620 47138
rect 434000 46818 434032 47054
rect 434268 46818 434352 47054
rect 434588 46818 434620 47054
rect 436560 47138 436622 47374
rect 436858 47138 436920 47374
rect 436560 47054 436920 47138
rect 436560 46818 436622 47054
rect 436858 46818 436920 47054
rect 409036 46786 409396 46818
rect 436560 46786 436920 46818
rect 535036 47374 535396 47406
rect 535036 47138 535098 47374
rect 535334 47138 535396 47374
rect 535036 47054 535396 47138
rect 535036 46818 535098 47054
rect 535334 46818 535396 47054
rect 542000 47138 542032 47374
rect 542268 47138 542352 47374
rect 542588 47138 542620 47374
rect 542000 47054 542620 47138
rect 542000 46818 542032 47054
rect 542268 46818 542352 47054
rect 542588 46818 542620 47054
rect 571500 47138 571532 47374
rect 571768 47138 571852 47374
rect 572088 47138 572120 47374
rect 571500 47054 572120 47138
rect 571500 46818 571532 47054
rect 571768 46818 571852 47054
rect 572088 46818 572120 47054
rect 535036 46786 535396 46818
rect 61280 43654 61640 43686
rect -2006 43418 -1974 43654
rect -1738 43418 -1654 43654
rect -1418 43418 -1386 43654
rect -2006 43334 -1386 43418
rect -2006 43098 -1974 43334
rect -1738 43098 -1654 43334
rect -1418 43098 -1386 43334
rect 9084 43418 9116 43654
rect 9352 43418 9436 43654
rect 9672 43418 9704 43654
rect 9084 43334 9704 43418
rect 9084 43098 9116 43334
rect 9352 43098 9436 43334
rect 9672 43098 9704 43334
rect 56620 43418 56652 43654
rect 56888 43418 56972 43654
rect 57208 43418 57240 43654
rect 56620 43334 57240 43418
rect 56620 43098 56652 43334
rect 56888 43098 56972 43334
rect 57208 43098 57240 43334
rect 61280 43418 61342 43654
rect 61578 43418 61640 43654
rect 61280 43334 61640 43418
rect 61280 43098 61342 43334
rect 61578 43098 61640 43334
rect -2006 3654 -1386 43098
rect 61280 43066 61640 43098
rect 158316 43654 158676 43686
rect 186280 43654 186640 43686
rect 158316 43418 158378 43654
rect 158614 43418 158676 43654
rect 158316 43334 158676 43418
rect 158316 43098 158378 43334
rect 158614 43098 158676 43334
rect 164620 43418 164652 43654
rect 164888 43418 164972 43654
rect 165208 43418 165240 43654
rect 164620 43334 165240 43418
rect 164620 43098 164652 43334
rect 164888 43098 164972 43334
rect 165208 43098 165240 43334
rect 186280 43418 186342 43654
rect 186578 43418 186640 43654
rect 186280 43334 186640 43418
rect 186280 43098 186342 43334
rect 186578 43098 186640 43334
rect 158316 43066 158676 43098
rect 186280 43066 186640 43098
rect 283316 43654 283676 43686
rect 311280 43654 311640 43686
rect 283316 43418 283378 43654
rect 283614 43418 283676 43654
rect 283316 43334 283676 43418
rect 283316 43098 283378 43334
rect 283614 43098 283676 43334
rect 308620 43418 308652 43654
rect 308888 43418 308972 43654
rect 309208 43418 309240 43654
rect 308620 43334 309240 43418
rect 308620 43098 308652 43334
rect 308888 43098 308972 43334
rect 309208 43098 309240 43334
rect 311280 43418 311342 43654
rect 311578 43418 311640 43654
rect 311280 43334 311640 43418
rect 311280 43098 311342 43334
rect 311578 43098 311640 43334
rect 283316 43066 283676 43098
rect 311280 43066 311640 43098
rect 408316 43654 408676 43686
rect 437280 43654 437640 43686
rect 408316 43418 408378 43654
rect 408614 43418 408676 43654
rect 408316 43334 408676 43418
rect 408316 43098 408378 43334
rect 408614 43098 408676 43334
rect 416620 43418 416652 43654
rect 416888 43418 416972 43654
rect 417208 43418 417240 43654
rect 416620 43334 417240 43418
rect 416620 43098 416652 43334
rect 416888 43098 416972 43334
rect 417208 43098 417240 43334
rect 437280 43418 437342 43654
rect 437578 43418 437640 43654
rect 437280 43334 437640 43418
rect 437280 43098 437342 43334
rect 437578 43098 437640 43334
rect 408316 43066 408676 43098
rect 437280 43066 437640 43098
rect 534316 43654 534676 43686
rect 534316 43418 534378 43654
rect 534614 43418 534676 43654
rect 534316 43334 534676 43418
rect 534316 43098 534378 43334
rect 534614 43098 534676 43334
rect 560620 43418 560652 43654
rect 560888 43418 560972 43654
rect 561208 43418 561240 43654
rect 560620 43334 561240 43418
rect 560620 43098 560652 43334
rect 560888 43098 560972 43334
rect 561208 43098 561240 43334
rect 570260 43418 570292 43654
rect 570528 43418 570612 43654
rect 570848 43418 570880 43654
rect 570260 43334 570880 43418
rect 570260 43098 570292 43334
rect 570528 43098 570612 43334
rect 570848 43098 570880 43334
rect 534316 43066 534676 43098
rect 580594 22254 581214 61698
rect 580594 22018 580626 22254
rect 580862 22018 580946 22254
rect 581182 22018 581214 22254
rect 580594 21934 581214 22018
rect 580594 21698 580626 21934
rect 580862 21698 580946 21934
rect 581182 21698 581214 21934
rect 61280 21244 61640 21300
rect 61280 21008 61342 21244
rect 61578 21008 61640 21244
rect 61280 20952 61640 21008
rect 62952 21244 63300 21300
rect 62952 21008 63008 21244
rect 63244 21008 63300 21244
rect 62952 20952 63300 21008
rect 187952 21244 188300 21300
rect 187952 21008 188008 21244
rect 188244 21008 188300 21244
rect 187952 20952 188300 21008
rect 311280 21244 311640 21300
rect 311280 21008 311342 21244
rect 311578 21008 311640 21244
rect 311280 20952 311640 21008
rect 312952 21244 313300 21300
rect 312952 21008 313008 21244
rect 313244 21008 313300 21244
rect 312952 20952 313300 21008
rect 438952 21244 439300 21300
rect 438952 21008 439008 21244
rect 439244 21008 439300 21244
rect 438952 20952 439300 21008
rect 62272 20564 62620 20620
rect 62272 20328 62328 20564
rect 62564 20328 62620 20564
rect 62272 20272 62620 20328
rect 185560 20564 185920 20620
rect 185560 20328 185622 20564
rect 185858 20328 185920 20564
rect 185560 20272 185920 20328
rect 187272 20564 187620 20620
rect 187272 20328 187328 20564
rect 187564 20328 187620 20564
rect 187272 20272 187620 20328
rect 312272 20564 312620 20620
rect 312272 20328 312328 20564
rect 312564 20328 312620 20564
rect 312272 20272 312620 20328
rect 436560 20564 436920 20620
rect 436560 20328 436622 20564
rect 436858 20328 436920 20564
rect 436560 20272 436920 20328
rect 438272 20564 438620 20620
rect 438272 20328 438328 20564
rect 438564 20328 438620 20564
rect 438272 20272 438620 20328
rect 62272 19834 62620 19858
rect 62272 19598 62328 19834
rect 62564 19598 62620 19834
rect 312272 19834 312620 19858
rect 62272 19574 62620 19598
rect 187952 19578 188300 19640
rect 187952 19342 188008 19578
rect 188244 19342 188300 19578
rect 312272 19598 312328 19834
rect 312564 19598 312620 19834
rect 312272 19574 312620 19598
rect 438952 19578 439300 19640
rect 187952 19280 188300 19342
rect 438952 19342 439008 19578
rect 439244 19342 439300 19578
rect 438952 19280 439300 19342
rect 9084 9444 9116 9680
rect 9352 9444 9436 9680
rect 9672 9444 9704 9680
rect 9084 9360 9704 9444
rect 9084 9124 9116 9360
rect 9352 9124 9436 9360
rect 9672 9124 9704 9360
rect 56620 9444 56652 9680
rect 56888 9444 56972 9680
rect 57208 9444 57240 9680
rect 56620 9360 57240 9444
rect 56620 9124 56652 9360
rect 56888 9124 56972 9360
rect 57208 9124 57240 9360
rect 92620 9444 92652 9680
rect 92888 9444 92972 9680
rect 93208 9444 93240 9680
rect 92620 9360 93240 9444
rect 92620 9124 92652 9360
rect 92888 9124 92972 9360
rect 93208 9124 93240 9360
rect 128620 9444 128652 9680
rect 128888 9444 128972 9680
rect 129208 9444 129240 9680
rect 128620 9360 129240 9444
rect 128620 9124 128652 9360
rect 128888 9124 128972 9360
rect 129208 9124 129240 9360
rect 164620 9444 164652 9680
rect 164888 9444 164972 9680
rect 165208 9444 165240 9680
rect 164620 9360 165240 9444
rect 164620 9124 164652 9360
rect 164888 9124 164972 9360
rect 165208 9124 165240 9360
rect 200620 9444 200652 9680
rect 200888 9444 200972 9680
rect 201208 9444 201240 9680
rect 200620 9360 201240 9444
rect 200620 9124 200652 9360
rect 200888 9124 200972 9360
rect 201208 9124 201240 9360
rect 236620 9444 236652 9680
rect 236888 9444 236972 9680
rect 237208 9444 237240 9680
rect 236620 9360 237240 9444
rect 236620 9124 236652 9360
rect 236888 9124 236972 9360
rect 237208 9124 237240 9360
rect 272620 9444 272652 9680
rect 272888 9444 272972 9680
rect 273208 9444 273240 9680
rect 272620 9360 273240 9444
rect 272620 9124 272652 9360
rect 272888 9124 272972 9360
rect 273208 9124 273240 9360
rect 308620 9444 308652 9680
rect 308888 9444 308972 9680
rect 309208 9444 309240 9680
rect 308620 9360 309240 9444
rect 308620 9124 308652 9360
rect 308888 9124 308972 9360
rect 309208 9124 309240 9360
rect 344620 9444 344652 9680
rect 344888 9444 344972 9680
rect 345208 9444 345240 9680
rect 344620 9360 345240 9444
rect 344620 9124 344652 9360
rect 344888 9124 344972 9360
rect 345208 9124 345240 9360
rect 380620 9444 380652 9680
rect 380888 9444 380972 9680
rect 381208 9444 381240 9680
rect 380620 9360 381240 9444
rect 380620 9124 380652 9360
rect 380888 9124 380972 9360
rect 381208 9124 381240 9360
rect 416620 9444 416652 9680
rect 416888 9444 416972 9680
rect 417208 9444 417240 9680
rect 416620 9360 417240 9444
rect 416620 9124 416652 9360
rect 416888 9124 416972 9360
rect 417208 9124 417240 9360
rect 452620 9444 452652 9680
rect 452888 9444 452972 9680
rect 453208 9444 453240 9680
rect 452620 9360 453240 9444
rect 452620 9124 452652 9360
rect 452888 9124 452972 9360
rect 453208 9124 453240 9360
rect 488620 9444 488652 9680
rect 488888 9444 488972 9680
rect 489208 9444 489240 9680
rect 488620 9360 489240 9444
rect 488620 9124 488652 9360
rect 488888 9124 488972 9360
rect 489208 9124 489240 9360
rect 524620 9444 524652 9680
rect 524888 9444 524972 9680
rect 525208 9444 525240 9680
rect 524620 9360 525240 9444
rect 524620 9124 524652 9360
rect 524888 9124 524972 9360
rect 525208 9124 525240 9360
rect 560620 9444 560652 9680
rect 560888 9444 560972 9680
rect 561208 9444 561240 9680
rect 560620 9360 561240 9444
rect 560620 9124 560652 9360
rect 560888 9124 560972 9360
rect 561208 9124 561240 9360
rect 570260 9444 570292 9680
rect 570528 9444 570612 9680
rect 570848 9444 570880 9680
rect 570260 9360 570880 9444
rect 570260 9124 570292 9360
rect 570528 9124 570612 9360
rect 570848 9124 570880 9360
rect 7844 8204 7876 8440
rect 8112 8204 8196 8440
rect 8432 8204 8464 8440
rect 7844 8120 8464 8204
rect 7844 7884 7876 8120
rect 8112 7884 8196 8120
rect 8432 7884 8464 8120
rect 38000 8204 38032 8440
rect 38268 8204 38352 8440
rect 38588 8204 38620 8440
rect 38000 8120 38620 8204
rect 38000 7884 38032 8120
rect 38268 7884 38352 8120
rect 38588 7884 38620 8120
rect 74000 8204 74032 8440
rect 74268 8204 74352 8440
rect 74588 8204 74620 8440
rect 74000 8120 74620 8204
rect 74000 7884 74032 8120
rect 74268 7884 74352 8120
rect 74588 7884 74620 8120
rect 110000 8204 110032 8440
rect 110268 8204 110352 8440
rect 110588 8204 110620 8440
rect 110000 8120 110620 8204
rect 110000 7884 110032 8120
rect 110268 7884 110352 8120
rect 110588 7884 110620 8120
rect 146000 8204 146032 8440
rect 146268 8204 146352 8440
rect 146588 8204 146620 8440
rect 146000 8120 146620 8204
rect 146000 7884 146032 8120
rect 146268 7884 146352 8120
rect 146588 7884 146620 8120
rect 182000 8204 182032 8440
rect 182268 8204 182352 8440
rect 182588 8204 182620 8440
rect 182000 8120 182620 8204
rect 182000 7884 182032 8120
rect 182268 7884 182352 8120
rect 182588 7884 182620 8120
rect 218000 8204 218032 8440
rect 218268 8204 218352 8440
rect 218588 8204 218620 8440
rect 218000 8120 218620 8204
rect 218000 7884 218032 8120
rect 218268 7884 218352 8120
rect 218588 7884 218620 8120
rect 254000 8204 254032 8440
rect 254268 8204 254352 8440
rect 254588 8204 254620 8440
rect 254000 8120 254620 8204
rect 254000 7884 254032 8120
rect 254268 7884 254352 8120
rect 254588 7884 254620 8120
rect 290000 8204 290032 8440
rect 290268 8204 290352 8440
rect 290588 8204 290620 8440
rect 290000 8120 290620 8204
rect 290000 7884 290032 8120
rect 290268 7884 290352 8120
rect 290588 7884 290620 8120
rect 326000 8204 326032 8440
rect 326268 8204 326352 8440
rect 326588 8204 326620 8440
rect 326000 8120 326620 8204
rect 326000 7884 326032 8120
rect 326268 7884 326352 8120
rect 326588 7884 326620 8120
rect 362000 8204 362032 8440
rect 362268 8204 362352 8440
rect 362588 8204 362620 8440
rect 362000 8120 362620 8204
rect 362000 7884 362032 8120
rect 362268 7884 362352 8120
rect 362588 7884 362620 8120
rect 398000 8204 398032 8440
rect 398268 8204 398352 8440
rect 398588 8204 398620 8440
rect 398000 8120 398620 8204
rect 398000 7884 398032 8120
rect 398268 7884 398352 8120
rect 398588 7884 398620 8120
rect 434000 8204 434032 8440
rect 434268 8204 434352 8440
rect 434588 8204 434620 8440
rect 434000 8120 434620 8204
rect 434000 7884 434032 8120
rect 434268 7884 434352 8120
rect 434588 7884 434620 8120
rect 470000 8204 470032 8440
rect 470268 8204 470352 8440
rect 470588 8204 470620 8440
rect 470000 8120 470620 8204
rect 470000 7884 470032 8120
rect 470268 7884 470352 8120
rect 470588 7884 470620 8120
rect 506000 8204 506032 8440
rect 506268 8204 506352 8440
rect 506588 8204 506620 8440
rect 506000 8120 506620 8204
rect 506000 7884 506032 8120
rect 506268 7884 506352 8120
rect 506588 7884 506620 8120
rect 542000 8204 542032 8440
rect 542268 8204 542352 8440
rect 542588 8204 542620 8440
rect 542000 8120 542620 8204
rect 542000 7884 542032 8120
rect 542268 7884 542352 8120
rect 542588 7884 542620 8120
rect 571500 8204 571532 8440
rect 571768 8204 571852 8440
rect 572088 8204 572120 8440
rect 571500 8120 572120 8204
rect 571500 7884 571532 8120
rect 571768 7884 571852 8120
rect 572088 7884 572120 8120
rect 7844 7138 7876 7374
rect 8112 7138 8196 7374
rect 8432 7138 8464 7374
rect 7844 7054 8464 7138
rect 7844 6818 7876 7054
rect 8112 6818 8196 7054
rect 8432 6818 8464 7054
rect 571500 7138 571532 7374
rect 571768 7138 571852 7374
rect 572088 7138 572120 7374
rect 571500 7054 572120 7138
rect 571500 6818 571532 7054
rect 571768 6818 571852 7054
rect 572088 6818 572120 7054
rect -2006 3418 -1974 3654
rect -1738 3418 -1654 3654
rect -1418 3418 -1386 3654
rect -2006 3334 -1386 3418
rect -2006 3098 -1974 3334
rect -1738 3098 -1654 3334
rect -1418 3098 -1386 3334
rect -2006 -346 -1386 3098
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect -5116 -3692 -5084 -3456
rect -4848 -3692 -4764 -3456
rect -4528 -3692 -4496 -3456
rect -5116 -3776 -4496 -3692
rect -5116 -4012 -5084 -3776
rect -4848 -4012 -4764 -3776
rect -4528 -4012 -4496 -3776
rect -5116 -4044 -4496 -4012
rect -8226 -6802 -8194 -6566
rect -7958 -6802 -7874 -6566
rect -7638 -6802 -7606 -6566
rect -8226 -6886 -7606 -6802
rect -8226 -7122 -8194 -6886
rect -7958 -7122 -7874 -6886
rect -7638 -7122 -7606 -6886
rect -8226 -7154 -7606 -7122
rect -11336 -9912 -11304 -9676
rect -11068 -9912 -10984 -9676
rect -10748 -9912 -10716 -9676
rect -11336 -9996 -10716 -9912
rect -11336 -10232 -11304 -9996
rect -11068 -10232 -10984 -9996
rect -10748 -10232 -10716 -9996
rect -11336 -10264 -10716 -10232
rect -14446 -13022 -14414 -12786
rect -14178 -13022 -14094 -12786
rect -13858 -13022 -13826 -12786
rect -14446 -13106 -13826 -13022
rect -14446 -13342 -14414 -13106
rect -14178 -13342 -14094 -13106
rect -13858 -13342 -13826 -13106
rect -14446 -13374 -13826 -13342
rect -17556 -16132 -17524 -15896
rect -17288 -16132 -17204 -15896
rect -16968 -16132 -16936 -15896
rect -17556 -16216 -16936 -16132
rect -17556 -16452 -17524 -16216
rect -17288 -16452 -17204 -16216
rect -16968 -16452 -16936 -16216
rect -17556 -16484 -16936 -16452
rect 580594 -15896 581214 21698
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 683654 585930 704282
rect 585310 683418 585342 683654
rect 585578 683418 585662 683654
rect 585898 683418 585930 683654
rect 585310 683334 585930 683418
rect 585310 683098 585342 683334
rect 585578 683098 585662 683334
rect 585898 683098 585930 683334
rect 585310 643654 585930 683098
rect 585310 643418 585342 643654
rect 585578 643418 585662 643654
rect 585898 643418 585930 643654
rect 585310 643334 585930 643418
rect 585310 643098 585342 643334
rect 585578 643098 585662 643334
rect 585898 643098 585930 643334
rect 585310 603654 585930 643098
rect 585310 603418 585342 603654
rect 585578 603418 585662 603654
rect 585898 603418 585930 603654
rect 585310 603334 585930 603418
rect 585310 603098 585342 603334
rect 585578 603098 585662 603334
rect 585898 603098 585930 603334
rect 585310 563654 585930 603098
rect 585310 563418 585342 563654
rect 585578 563418 585662 563654
rect 585898 563418 585930 563654
rect 585310 563334 585930 563418
rect 585310 563098 585342 563334
rect 585578 563098 585662 563334
rect 585898 563098 585930 563334
rect 585310 523654 585930 563098
rect 585310 523418 585342 523654
rect 585578 523418 585662 523654
rect 585898 523418 585930 523654
rect 585310 523334 585930 523418
rect 585310 523098 585342 523334
rect 585578 523098 585662 523334
rect 585898 523098 585930 523334
rect 585310 483654 585930 523098
rect 585310 483418 585342 483654
rect 585578 483418 585662 483654
rect 585898 483418 585930 483654
rect 585310 483334 585930 483418
rect 585310 483098 585342 483334
rect 585578 483098 585662 483334
rect 585898 483098 585930 483334
rect 585310 443654 585930 483098
rect 585310 443418 585342 443654
rect 585578 443418 585662 443654
rect 585898 443418 585930 443654
rect 585310 443334 585930 443418
rect 585310 443098 585342 443334
rect 585578 443098 585662 443334
rect 585898 443098 585930 443334
rect 585310 403654 585930 443098
rect 585310 403418 585342 403654
rect 585578 403418 585662 403654
rect 585898 403418 585930 403654
rect 585310 403334 585930 403418
rect 585310 403098 585342 403334
rect 585578 403098 585662 403334
rect 585898 403098 585930 403334
rect 585310 363654 585930 403098
rect 585310 363418 585342 363654
rect 585578 363418 585662 363654
rect 585898 363418 585930 363654
rect 585310 363334 585930 363418
rect 585310 363098 585342 363334
rect 585578 363098 585662 363334
rect 585898 363098 585930 363334
rect 585310 323654 585930 363098
rect 585310 323418 585342 323654
rect 585578 323418 585662 323654
rect 585898 323418 585930 323654
rect 585310 323334 585930 323418
rect 585310 323098 585342 323334
rect 585578 323098 585662 323334
rect 585898 323098 585930 323334
rect 585310 283654 585930 323098
rect 585310 283418 585342 283654
rect 585578 283418 585662 283654
rect 585898 283418 585930 283654
rect 585310 283334 585930 283418
rect 585310 283098 585342 283334
rect 585578 283098 585662 283334
rect 585898 283098 585930 283334
rect 585310 243654 585930 283098
rect 585310 243418 585342 243654
rect 585578 243418 585662 243654
rect 585898 243418 585930 243654
rect 585310 243334 585930 243418
rect 585310 243098 585342 243334
rect 585578 243098 585662 243334
rect 585898 243098 585930 243334
rect 585310 203654 585930 243098
rect 585310 203418 585342 203654
rect 585578 203418 585662 203654
rect 585898 203418 585930 203654
rect 585310 203334 585930 203418
rect 585310 203098 585342 203334
rect 585578 203098 585662 203334
rect 585898 203098 585930 203334
rect 585310 163654 585930 203098
rect 585310 163418 585342 163654
rect 585578 163418 585662 163654
rect 585898 163418 585930 163654
rect 585310 163334 585930 163418
rect 585310 163098 585342 163334
rect 585578 163098 585662 163334
rect 585898 163098 585930 163334
rect 585310 123654 585930 163098
rect 585310 123418 585342 123654
rect 585578 123418 585662 123654
rect 585898 123418 585930 123654
rect 585310 123334 585930 123418
rect 585310 123098 585342 123334
rect 585578 123098 585662 123334
rect 585898 123098 585930 123334
rect 585310 83654 585930 123098
rect 585310 83418 585342 83654
rect 585578 83418 585662 83654
rect 585898 83418 585930 83654
rect 585310 83334 585930 83418
rect 585310 83098 585342 83334
rect 585578 83098 585662 83334
rect 585898 83098 585930 83334
rect 585310 43654 585930 83098
rect 585310 43418 585342 43654
rect 585578 43418 585662 43654
rect 585898 43418 585930 43654
rect 585310 43334 585930 43418
rect 585310 43098 585342 43334
rect 585578 43098 585662 43334
rect 585898 43098 585930 43334
rect 585310 3654 585930 43098
rect 585310 3418 585342 3654
rect 585578 3418 585662 3654
rect 585898 3418 585930 3654
rect 585310 3334 585930 3418
rect 585310 3098 585342 3334
rect 585578 3098 585662 3334
rect 585898 3098 585930 3334
rect 585310 -346 585930 3098
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 588420 687374 589040 707392
rect 588420 687138 588452 687374
rect 588688 687138 588772 687374
rect 589008 687138 589040 687374
rect 588420 687054 589040 687138
rect 588420 686818 588452 687054
rect 588688 686818 588772 687054
rect 589008 686818 589040 687054
rect 588420 647374 589040 686818
rect 588420 647138 588452 647374
rect 588688 647138 588772 647374
rect 589008 647138 589040 647374
rect 588420 647054 589040 647138
rect 588420 646818 588452 647054
rect 588688 646818 588772 647054
rect 589008 646818 589040 647054
rect 588420 607374 589040 646818
rect 588420 607138 588452 607374
rect 588688 607138 588772 607374
rect 589008 607138 589040 607374
rect 588420 607054 589040 607138
rect 588420 606818 588452 607054
rect 588688 606818 588772 607054
rect 589008 606818 589040 607054
rect 588420 567374 589040 606818
rect 588420 567138 588452 567374
rect 588688 567138 588772 567374
rect 589008 567138 589040 567374
rect 588420 567054 589040 567138
rect 588420 566818 588452 567054
rect 588688 566818 588772 567054
rect 589008 566818 589040 567054
rect 588420 527374 589040 566818
rect 588420 527138 588452 527374
rect 588688 527138 588772 527374
rect 589008 527138 589040 527374
rect 588420 527054 589040 527138
rect 588420 526818 588452 527054
rect 588688 526818 588772 527054
rect 589008 526818 589040 527054
rect 588420 487374 589040 526818
rect 588420 487138 588452 487374
rect 588688 487138 588772 487374
rect 589008 487138 589040 487374
rect 588420 487054 589040 487138
rect 588420 486818 588452 487054
rect 588688 486818 588772 487054
rect 589008 486818 589040 487054
rect 588420 447374 589040 486818
rect 588420 447138 588452 447374
rect 588688 447138 588772 447374
rect 589008 447138 589040 447374
rect 588420 447054 589040 447138
rect 588420 446818 588452 447054
rect 588688 446818 588772 447054
rect 589008 446818 589040 447054
rect 588420 407374 589040 446818
rect 588420 407138 588452 407374
rect 588688 407138 588772 407374
rect 589008 407138 589040 407374
rect 588420 407054 589040 407138
rect 588420 406818 588452 407054
rect 588688 406818 588772 407054
rect 589008 406818 589040 407054
rect 588420 367374 589040 406818
rect 588420 367138 588452 367374
rect 588688 367138 588772 367374
rect 589008 367138 589040 367374
rect 588420 367054 589040 367138
rect 588420 366818 588452 367054
rect 588688 366818 588772 367054
rect 589008 366818 589040 367054
rect 588420 327374 589040 366818
rect 588420 327138 588452 327374
rect 588688 327138 588772 327374
rect 589008 327138 589040 327374
rect 588420 327054 589040 327138
rect 588420 326818 588452 327054
rect 588688 326818 588772 327054
rect 589008 326818 589040 327054
rect 588420 287374 589040 326818
rect 588420 287138 588452 287374
rect 588688 287138 588772 287374
rect 589008 287138 589040 287374
rect 588420 287054 589040 287138
rect 588420 286818 588452 287054
rect 588688 286818 588772 287054
rect 589008 286818 589040 287054
rect 588420 247374 589040 286818
rect 588420 247138 588452 247374
rect 588688 247138 588772 247374
rect 589008 247138 589040 247374
rect 588420 247054 589040 247138
rect 588420 246818 588452 247054
rect 588688 246818 588772 247054
rect 589008 246818 589040 247054
rect 588420 207374 589040 246818
rect 588420 207138 588452 207374
rect 588688 207138 588772 207374
rect 589008 207138 589040 207374
rect 588420 207054 589040 207138
rect 588420 206818 588452 207054
rect 588688 206818 588772 207054
rect 589008 206818 589040 207054
rect 588420 167374 589040 206818
rect 588420 167138 588452 167374
rect 588688 167138 588772 167374
rect 589008 167138 589040 167374
rect 588420 167054 589040 167138
rect 588420 166818 588452 167054
rect 588688 166818 588772 167054
rect 589008 166818 589040 167054
rect 588420 127374 589040 166818
rect 588420 127138 588452 127374
rect 588688 127138 588772 127374
rect 589008 127138 589040 127374
rect 588420 127054 589040 127138
rect 588420 126818 588452 127054
rect 588688 126818 588772 127054
rect 589008 126818 589040 127054
rect 588420 87374 589040 126818
rect 588420 87138 588452 87374
rect 588688 87138 588772 87374
rect 589008 87138 589040 87374
rect 588420 87054 589040 87138
rect 588420 86818 588452 87054
rect 588688 86818 588772 87054
rect 589008 86818 589040 87054
rect 588420 47374 589040 86818
rect 588420 47138 588452 47374
rect 588688 47138 588772 47374
rect 589008 47138 589040 47374
rect 588420 47054 589040 47138
rect 588420 46818 588452 47054
rect 588688 46818 588772 47054
rect 589008 46818 589040 47054
rect 588420 7374 589040 46818
rect 588420 7138 588452 7374
rect 588688 7138 588772 7374
rect 589008 7138 589040 7374
rect 588420 7054 589040 7138
rect 588420 6818 588452 7054
rect 588688 6818 588772 7054
rect 589008 6818 589040 7054
rect 588420 -3456 589040 6818
rect 588420 -3692 588452 -3456
rect 588688 -3692 588772 -3456
rect 589008 -3692 589040 -3456
rect 588420 -3776 589040 -3692
rect 588420 -4012 588452 -3776
rect 588688 -4012 588772 -3776
rect 589008 -4012 589040 -3776
rect 588420 -4044 589040 -4012
rect 591530 691094 592150 710502
rect 591530 690858 591562 691094
rect 591798 690858 591882 691094
rect 592118 690858 592150 691094
rect 591530 690774 592150 690858
rect 591530 690538 591562 690774
rect 591798 690538 591882 690774
rect 592118 690538 592150 690774
rect 591530 651094 592150 690538
rect 591530 650858 591562 651094
rect 591798 650858 591882 651094
rect 592118 650858 592150 651094
rect 591530 650774 592150 650858
rect 591530 650538 591562 650774
rect 591798 650538 591882 650774
rect 592118 650538 592150 650774
rect 591530 611094 592150 650538
rect 591530 610858 591562 611094
rect 591798 610858 591882 611094
rect 592118 610858 592150 611094
rect 591530 610774 592150 610858
rect 591530 610538 591562 610774
rect 591798 610538 591882 610774
rect 592118 610538 592150 610774
rect 591530 571094 592150 610538
rect 591530 570858 591562 571094
rect 591798 570858 591882 571094
rect 592118 570858 592150 571094
rect 591530 570774 592150 570858
rect 591530 570538 591562 570774
rect 591798 570538 591882 570774
rect 592118 570538 592150 570774
rect 591530 531094 592150 570538
rect 591530 530858 591562 531094
rect 591798 530858 591882 531094
rect 592118 530858 592150 531094
rect 591530 530774 592150 530858
rect 591530 530538 591562 530774
rect 591798 530538 591882 530774
rect 592118 530538 592150 530774
rect 591530 491094 592150 530538
rect 591530 490858 591562 491094
rect 591798 490858 591882 491094
rect 592118 490858 592150 491094
rect 591530 490774 592150 490858
rect 591530 490538 591562 490774
rect 591798 490538 591882 490774
rect 592118 490538 592150 490774
rect 591530 451094 592150 490538
rect 591530 450858 591562 451094
rect 591798 450858 591882 451094
rect 592118 450858 592150 451094
rect 591530 450774 592150 450858
rect 591530 450538 591562 450774
rect 591798 450538 591882 450774
rect 592118 450538 592150 450774
rect 591530 411094 592150 450538
rect 591530 410858 591562 411094
rect 591798 410858 591882 411094
rect 592118 410858 592150 411094
rect 591530 410774 592150 410858
rect 591530 410538 591562 410774
rect 591798 410538 591882 410774
rect 592118 410538 592150 410774
rect 591530 371094 592150 410538
rect 591530 370858 591562 371094
rect 591798 370858 591882 371094
rect 592118 370858 592150 371094
rect 591530 370774 592150 370858
rect 591530 370538 591562 370774
rect 591798 370538 591882 370774
rect 592118 370538 592150 370774
rect 591530 331094 592150 370538
rect 591530 330858 591562 331094
rect 591798 330858 591882 331094
rect 592118 330858 592150 331094
rect 591530 330774 592150 330858
rect 591530 330538 591562 330774
rect 591798 330538 591882 330774
rect 592118 330538 592150 330774
rect 591530 291094 592150 330538
rect 591530 290858 591562 291094
rect 591798 290858 591882 291094
rect 592118 290858 592150 291094
rect 591530 290774 592150 290858
rect 591530 290538 591562 290774
rect 591798 290538 591882 290774
rect 592118 290538 592150 290774
rect 591530 251094 592150 290538
rect 591530 250858 591562 251094
rect 591798 250858 591882 251094
rect 592118 250858 592150 251094
rect 591530 250774 592150 250858
rect 591530 250538 591562 250774
rect 591798 250538 591882 250774
rect 592118 250538 592150 250774
rect 591530 211094 592150 250538
rect 591530 210858 591562 211094
rect 591798 210858 591882 211094
rect 592118 210858 592150 211094
rect 591530 210774 592150 210858
rect 591530 210538 591562 210774
rect 591798 210538 591882 210774
rect 592118 210538 592150 210774
rect 591530 171094 592150 210538
rect 591530 170858 591562 171094
rect 591798 170858 591882 171094
rect 592118 170858 592150 171094
rect 591530 170774 592150 170858
rect 591530 170538 591562 170774
rect 591798 170538 591882 170774
rect 592118 170538 592150 170774
rect 591530 131094 592150 170538
rect 591530 130858 591562 131094
rect 591798 130858 591882 131094
rect 592118 130858 592150 131094
rect 591530 130774 592150 130858
rect 591530 130538 591562 130774
rect 591798 130538 591882 130774
rect 592118 130538 592150 130774
rect 591530 91094 592150 130538
rect 591530 90858 591562 91094
rect 591798 90858 591882 91094
rect 592118 90858 592150 91094
rect 591530 90774 592150 90858
rect 591530 90538 591562 90774
rect 591798 90538 591882 90774
rect 592118 90538 592150 90774
rect 591530 51094 592150 90538
rect 591530 50858 591562 51094
rect 591798 50858 591882 51094
rect 592118 50858 592150 51094
rect 591530 50774 592150 50858
rect 591530 50538 591562 50774
rect 591798 50538 591882 50774
rect 592118 50538 592150 50774
rect 591530 11094 592150 50538
rect 591530 10858 591562 11094
rect 591798 10858 591882 11094
rect 592118 10858 592150 11094
rect 591530 10774 592150 10858
rect 591530 10538 591562 10774
rect 591798 10538 591882 10774
rect 592118 10538 592150 10774
rect 591530 -6566 592150 10538
rect 591530 -6802 591562 -6566
rect 591798 -6802 591882 -6566
rect 592118 -6802 592150 -6566
rect 591530 -6886 592150 -6802
rect 591530 -7122 591562 -6886
rect 591798 -7122 591882 -6886
rect 592118 -7122 592150 -6886
rect 591530 -7154 592150 -7122
rect 594640 694814 595260 713612
rect 594640 694578 594672 694814
rect 594908 694578 594992 694814
rect 595228 694578 595260 694814
rect 594640 694494 595260 694578
rect 594640 694258 594672 694494
rect 594908 694258 594992 694494
rect 595228 694258 595260 694494
rect 594640 654814 595260 694258
rect 594640 654578 594672 654814
rect 594908 654578 594992 654814
rect 595228 654578 595260 654814
rect 594640 654494 595260 654578
rect 594640 654258 594672 654494
rect 594908 654258 594992 654494
rect 595228 654258 595260 654494
rect 594640 614814 595260 654258
rect 594640 614578 594672 614814
rect 594908 614578 594992 614814
rect 595228 614578 595260 614814
rect 594640 614494 595260 614578
rect 594640 614258 594672 614494
rect 594908 614258 594992 614494
rect 595228 614258 595260 614494
rect 594640 574814 595260 614258
rect 594640 574578 594672 574814
rect 594908 574578 594992 574814
rect 595228 574578 595260 574814
rect 594640 574494 595260 574578
rect 594640 574258 594672 574494
rect 594908 574258 594992 574494
rect 595228 574258 595260 574494
rect 594640 534814 595260 574258
rect 594640 534578 594672 534814
rect 594908 534578 594992 534814
rect 595228 534578 595260 534814
rect 594640 534494 595260 534578
rect 594640 534258 594672 534494
rect 594908 534258 594992 534494
rect 595228 534258 595260 534494
rect 594640 494814 595260 534258
rect 594640 494578 594672 494814
rect 594908 494578 594992 494814
rect 595228 494578 595260 494814
rect 594640 494494 595260 494578
rect 594640 494258 594672 494494
rect 594908 494258 594992 494494
rect 595228 494258 595260 494494
rect 594640 454814 595260 494258
rect 594640 454578 594672 454814
rect 594908 454578 594992 454814
rect 595228 454578 595260 454814
rect 594640 454494 595260 454578
rect 594640 454258 594672 454494
rect 594908 454258 594992 454494
rect 595228 454258 595260 454494
rect 594640 414814 595260 454258
rect 594640 414578 594672 414814
rect 594908 414578 594992 414814
rect 595228 414578 595260 414814
rect 594640 414494 595260 414578
rect 594640 414258 594672 414494
rect 594908 414258 594992 414494
rect 595228 414258 595260 414494
rect 594640 374814 595260 414258
rect 594640 374578 594672 374814
rect 594908 374578 594992 374814
rect 595228 374578 595260 374814
rect 594640 374494 595260 374578
rect 594640 374258 594672 374494
rect 594908 374258 594992 374494
rect 595228 374258 595260 374494
rect 594640 334814 595260 374258
rect 594640 334578 594672 334814
rect 594908 334578 594992 334814
rect 595228 334578 595260 334814
rect 594640 334494 595260 334578
rect 594640 334258 594672 334494
rect 594908 334258 594992 334494
rect 595228 334258 595260 334494
rect 594640 294814 595260 334258
rect 594640 294578 594672 294814
rect 594908 294578 594992 294814
rect 595228 294578 595260 294814
rect 594640 294494 595260 294578
rect 594640 294258 594672 294494
rect 594908 294258 594992 294494
rect 595228 294258 595260 294494
rect 594640 254814 595260 294258
rect 594640 254578 594672 254814
rect 594908 254578 594992 254814
rect 595228 254578 595260 254814
rect 594640 254494 595260 254578
rect 594640 254258 594672 254494
rect 594908 254258 594992 254494
rect 595228 254258 595260 254494
rect 594640 214814 595260 254258
rect 594640 214578 594672 214814
rect 594908 214578 594992 214814
rect 595228 214578 595260 214814
rect 594640 214494 595260 214578
rect 594640 214258 594672 214494
rect 594908 214258 594992 214494
rect 595228 214258 595260 214494
rect 594640 174814 595260 214258
rect 594640 174578 594672 174814
rect 594908 174578 594992 174814
rect 595228 174578 595260 174814
rect 594640 174494 595260 174578
rect 594640 174258 594672 174494
rect 594908 174258 594992 174494
rect 595228 174258 595260 174494
rect 594640 134814 595260 174258
rect 594640 134578 594672 134814
rect 594908 134578 594992 134814
rect 595228 134578 595260 134814
rect 594640 134494 595260 134578
rect 594640 134258 594672 134494
rect 594908 134258 594992 134494
rect 595228 134258 595260 134494
rect 594640 94814 595260 134258
rect 594640 94578 594672 94814
rect 594908 94578 594992 94814
rect 595228 94578 595260 94814
rect 594640 94494 595260 94578
rect 594640 94258 594672 94494
rect 594908 94258 594992 94494
rect 595228 94258 595260 94494
rect 594640 54814 595260 94258
rect 594640 54578 594672 54814
rect 594908 54578 594992 54814
rect 595228 54578 595260 54814
rect 594640 54494 595260 54578
rect 594640 54258 594672 54494
rect 594908 54258 594992 54494
rect 595228 54258 595260 54494
rect 594640 14814 595260 54258
rect 594640 14578 594672 14814
rect 594908 14578 594992 14814
rect 595228 14578 595260 14814
rect 594640 14494 595260 14578
rect 594640 14258 594672 14494
rect 594908 14258 594992 14494
rect 595228 14258 595260 14494
rect 594640 -9676 595260 14258
rect 594640 -9912 594672 -9676
rect 594908 -9912 594992 -9676
rect 595228 -9912 595260 -9676
rect 594640 -9996 595260 -9912
rect 594640 -10232 594672 -9996
rect 594908 -10232 594992 -9996
rect 595228 -10232 595260 -9996
rect 594640 -10264 595260 -10232
rect 597750 698534 598370 716722
rect 597750 698298 597782 698534
rect 598018 698298 598102 698534
rect 598338 698298 598370 698534
rect 597750 698214 598370 698298
rect 597750 697978 597782 698214
rect 598018 697978 598102 698214
rect 598338 697978 598370 698214
rect 597750 658534 598370 697978
rect 597750 658298 597782 658534
rect 598018 658298 598102 658534
rect 598338 658298 598370 658534
rect 597750 658214 598370 658298
rect 597750 657978 597782 658214
rect 598018 657978 598102 658214
rect 598338 657978 598370 658214
rect 597750 618534 598370 657978
rect 597750 618298 597782 618534
rect 598018 618298 598102 618534
rect 598338 618298 598370 618534
rect 597750 618214 598370 618298
rect 597750 617978 597782 618214
rect 598018 617978 598102 618214
rect 598338 617978 598370 618214
rect 597750 578534 598370 617978
rect 597750 578298 597782 578534
rect 598018 578298 598102 578534
rect 598338 578298 598370 578534
rect 597750 578214 598370 578298
rect 597750 577978 597782 578214
rect 598018 577978 598102 578214
rect 598338 577978 598370 578214
rect 597750 538534 598370 577978
rect 597750 538298 597782 538534
rect 598018 538298 598102 538534
rect 598338 538298 598370 538534
rect 597750 538214 598370 538298
rect 597750 537978 597782 538214
rect 598018 537978 598102 538214
rect 598338 537978 598370 538214
rect 597750 498534 598370 537978
rect 597750 498298 597782 498534
rect 598018 498298 598102 498534
rect 598338 498298 598370 498534
rect 597750 498214 598370 498298
rect 597750 497978 597782 498214
rect 598018 497978 598102 498214
rect 598338 497978 598370 498214
rect 597750 458534 598370 497978
rect 597750 458298 597782 458534
rect 598018 458298 598102 458534
rect 598338 458298 598370 458534
rect 597750 458214 598370 458298
rect 597750 457978 597782 458214
rect 598018 457978 598102 458214
rect 598338 457978 598370 458214
rect 597750 418534 598370 457978
rect 597750 418298 597782 418534
rect 598018 418298 598102 418534
rect 598338 418298 598370 418534
rect 597750 418214 598370 418298
rect 597750 417978 597782 418214
rect 598018 417978 598102 418214
rect 598338 417978 598370 418214
rect 597750 378534 598370 417978
rect 597750 378298 597782 378534
rect 598018 378298 598102 378534
rect 598338 378298 598370 378534
rect 597750 378214 598370 378298
rect 597750 377978 597782 378214
rect 598018 377978 598102 378214
rect 598338 377978 598370 378214
rect 597750 338534 598370 377978
rect 597750 338298 597782 338534
rect 598018 338298 598102 338534
rect 598338 338298 598370 338534
rect 597750 338214 598370 338298
rect 597750 337978 597782 338214
rect 598018 337978 598102 338214
rect 598338 337978 598370 338214
rect 597750 298534 598370 337978
rect 597750 298298 597782 298534
rect 598018 298298 598102 298534
rect 598338 298298 598370 298534
rect 597750 298214 598370 298298
rect 597750 297978 597782 298214
rect 598018 297978 598102 298214
rect 598338 297978 598370 298214
rect 597750 258534 598370 297978
rect 597750 258298 597782 258534
rect 598018 258298 598102 258534
rect 598338 258298 598370 258534
rect 597750 258214 598370 258298
rect 597750 257978 597782 258214
rect 598018 257978 598102 258214
rect 598338 257978 598370 258214
rect 597750 218534 598370 257978
rect 597750 218298 597782 218534
rect 598018 218298 598102 218534
rect 598338 218298 598370 218534
rect 597750 218214 598370 218298
rect 597750 217978 597782 218214
rect 598018 217978 598102 218214
rect 598338 217978 598370 218214
rect 597750 178534 598370 217978
rect 597750 178298 597782 178534
rect 598018 178298 598102 178534
rect 598338 178298 598370 178534
rect 597750 178214 598370 178298
rect 597750 177978 597782 178214
rect 598018 177978 598102 178214
rect 598338 177978 598370 178214
rect 597750 138534 598370 177978
rect 597750 138298 597782 138534
rect 598018 138298 598102 138534
rect 598338 138298 598370 138534
rect 597750 138214 598370 138298
rect 597750 137978 597782 138214
rect 598018 137978 598102 138214
rect 598338 137978 598370 138214
rect 597750 98534 598370 137978
rect 597750 98298 597782 98534
rect 598018 98298 598102 98534
rect 598338 98298 598370 98534
rect 597750 98214 598370 98298
rect 597750 97978 597782 98214
rect 598018 97978 598102 98214
rect 598338 97978 598370 98214
rect 597750 58534 598370 97978
rect 597750 58298 597782 58534
rect 598018 58298 598102 58534
rect 598338 58298 598370 58534
rect 597750 58214 598370 58298
rect 597750 57978 597782 58214
rect 598018 57978 598102 58214
rect 598338 57978 598370 58214
rect 597750 18534 598370 57978
rect 597750 18298 597782 18534
rect 598018 18298 598102 18534
rect 598338 18298 598370 18534
rect 597750 18214 598370 18298
rect 597750 17978 597782 18214
rect 598018 17978 598102 18214
rect 598338 17978 598370 18214
rect 597750 -12786 598370 17978
rect 597750 -13022 597782 -12786
rect 598018 -13022 598102 -12786
rect 598338 -13022 598370 -12786
rect 597750 -13106 598370 -13022
rect 597750 -13342 597782 -13106
rect 598018 -13342 598102 -13106
rect 598338 -13342 598370 -13106
rect 597750 -13374 598370 -13342
rect 600860 662254 601480 719832
rect 600860 662018 600892 662254
rect 601128 662018 601212 662254
rect 601448 662018 601480 662254
rect 600860 661934 601480 662018
rect 600860 661698 600892 661934
rect 601128 661698 601212 661934
rect 601448 661698 601480 661934
rect 600860 622254 601480 661698
rect 600860 622018 600892 622254
rect 601128 622018 601212 622254
rect 601448 622018 601480 622254
rect 600860 621934 601480 622018
rect 600860 621698 600892 621934
rect 601128 621698 601212 621934
rect 601448 621698 601480 621934
rect 600860 582254 601480 621698
rect 600860 582018 600892 582254
rect 601128 582018 601212 582254
rect 601448 582018 601480 582254
rect 600860 581934 601480 582018
rect 600860 581698 600892 581934
rect 601128 581698 601212 581934
rect 601448 581698 601480 581934
rect 600860 542254 601480 581698
rect 600860 542018 600892 542254
rect 601128 542018 601212 542254
rect 601448 542018 601480 542254
rect 600860 541934 601480 542018
rect 600860 541698 600892 541934
rect 601128 541698 601212 541934
rect 601448 541698 601480 541934
rect 600860 502254 601480 541698
rect 600860 502018 600892 502254
rect 601128 502018 601212 502254
rect 601448 502018 601480 502254
rect 600860 501934 601480 502018
rect 600860 501698 600892 501934
rect 601128 501698 601212 501934
rect 601448 501698 601480 501934
rect 600860 462254 601480 501698
rect 600860 462018 600892 462254
rect 601128 462018 601212 462254
rect 601448 462018 601480 462254
rect 600860 461934 601480 462018
rect 600860 461698 600892 461934
rect 601128 461698 601212 461934
rect 601448 461698 601480 461934
rect 600860 422254 601480 461698
rect 600860 422018 600892 422254
rect 601128 422018 601212 422254
rect 601448 422018 601480 422254
rect 600860 421934 601480 422018
rect 600860 421698 600892 421934
rect 601128 421698 601212 421934
rect 601448 421698 601480 421934
rect 600860 382254 601480 421698
rect 600860 382018 600892 382254
rect 601128 382018 601212 382254
rect 601448 382018 601480 382254
rect 600860 381934 601480 382018
rect 600860 381698 600892 381934
rect 601128 381698 601212 381934
rect 601448 381698 601480 381934
rect 600860 342254 601480 381698
rect 600860 342018 600892 342254
rect 601128 342018 601212 342254
rect 601448 342018 601480 342254
rect 600860 341934 601480 342018
rect 600860 341698 600892 341934
rect 601128 341698 601212 341934
rect 601448 341698 601480 341934
rect 600860 302254 601480 341698
rect 600860 302018 600892 302254
rect 601128 302018 601212 302254
rect 601448 302018 601480 302254
rect 600860 301934 601480 302018
rect 600860 301698 600892 301934
rect 601128 301698 601212 301934
rect 601448 301698 601480 301934
rect 600860 262254 601480 301698
rect 600860 262018 600892 262254
rect 601128 262018 601212 262254
rect 601448 262018 601480 262254
rect 600860 261934 601480 262018
rect 600860 261698 600892 261934
rect 601128 261698 601212 261934
rect 601448 261698 601480 261934
rect 600860 222254 601480 261698
rect 600860 222018 600892 222254
rect 601128 222018 601212 222254
rect 601448 222018 601480 222254
rect 600860 221934 601480 222018
rect 600860 221698 600892 221934
rect 601128 221698 601212 221934
rect 601448 221698 601480 221934
rect 600860 182254 601480 221698
rect 600860 182018 600892 182254
rect 601128 182018 601212 182254
rect 601448 182018 601480 182254
rect 600860 181934 601480 182018
rect 600860 181698 600892 181934
rect 601128 181698 601212 181934
rect 601448 181698 601480 181934
rect 600860 142254 601480 181698
rect 600860 142018 600892 142254
rect 601128 142018 601212 142254
rect 601448 142018 601480 142254
rect 600860 141934 601480 142018
rect 600860 141698 600892 141934
rect 601128 141698 601212 141934
rect 601448 141698 601480 141934
rect 600860 102254 601480 141698
rect 600860 102018 600892 102254
rect 601128 102018 601212 102254
rect 601448 102018 601480 102254
rect 600860 101934 601480 102018
rect 600860 101698 600892 101934
rect 601128 101698 601212 101934
rect 601448 101698 601480 101934
rect 600860 62254 601480 101698
rect 600860 62018 600892 62254
rect 601128 62018 601212 62254
rect 601448 62018 601480 62254
rect 600860 61934 601480 62018
rect 600860 61698 600892 61934
rect 601128 61698 601212 61934
rect 601448 61698 601480 61934
rect 600860 22254 601480 61698
rect 600860 22018 600892 22254
rect 601128 22018 601212 22254
rect 601448 22018 601480 22254
rect 600860 21934 601480 22018
rect 600860 21698 600892 21934
rect 601128 21698 601212 21934
rect 601448 21698 601480 21934
rect 580594 -16132 580626 -15896
rect 580862 -16132 580946 -15896
rect 581182 -16132 581214 -15896
rect 580594 -16216 581214 -16132
rect 580594 -16452 580626 -16216
rect 580862 -16452 580946 -16216
rect 581182 -16452 581214 -16216
rect -20666 -19242 -20634 -19006
rect -20398 -19242 -20314 -19006
rect -20078 -19242 -20046 -19006
rect -20666 -19326 -20046 -19242
rect -20666 -19562 -20634 -19326
rect -20398 -19562 -20314 -19326
rect -20078 -19562 -20046 -19326
rect -20666 -19594 -20046 -19562
rect -23776 -22352 -23744 -22116
rect -23508 -22352 -23424 -22116
rect -23188 -22352 -23156 -22116
rect -23776 -22436 -23156 -22352
rect -23776 -22672 -23744 -22436
rect -23508 -22672 -23424 -22436
rect -23188 -22672 -23156 -22436
rect -23776 -22704 -23156 -22672
rect 580594 -22704 581214 -16452
rect 600860 -15896 601480 21698
rect 600860 -16132 600892 -15896
rect 601128 -16132 601212 -15896
rect 601448 -16132 601480 -15896
rect 600860 -16216 601480 -16132
rect 600860 -16452 600892 -16216
rect 601128 -16452 601212 -16216
rect 601448 -16452 601480 -16216
rect 600860 -16484 601480 -16452
rect 603970 665974 604590 722942
rect 603970 665738 604002 665974
rect 604238 665738 604322 665974
rect 604558 665738 604590 665974
rect 603970 665654 604590 665738
rect 603970 665418 604002 665654
rect 604238 665418 604322 665654
rect 604558 665418 604590 665654
rect 603970 625974 604590 665418
rect 603970 625738 604002 625974
rect 604238 625738 604322 625974
rect 604558 625738 604590 625974
rect 603970 625654 604590 625738
rect 603970 625418 604002 625654
rect 604238 625418 604322 625654
rect 604558 625418 604590 625654
rect 603970 585974 604590 625418
rect 603970 585738 604002 585974
rect 604238 585738 604322 585974
rect 604558 585738 604590 585974
rect 603970 585654 604590 585738
rect 603970 585418 604002 585654
rect 604238 585418 604322 585654
rect 604558 585418 604590 585654
rect 603970 545974 604590 585418
rect 603970 545738 604002 545974
rect 604238 545738 604322 545974
rect 604558 545738 604590 545974
rect 603970 545654 604590 545738
rect 603970 545418 604002 545654
rect 604238 545418 604322 545654
rect 604558 545418 604590 545654
rect 603970 505974 604590 545418
rect 603970 505738 604002 505974
rect 604238 505738 604322 505974
rect 604558 505738 604590 505974
rect 603970 505654 604590 505738
rect 603970 505418 604002 505654
rect 604238 505418 604322 505654
rect 604558 505418 604590 505654
rect 603970 465974 604590 505418
rect 603970 465738 604002 465974
rect 604238 465738 604322 465974
rect 604558 465738 604590 465974
rect 603970 465654 604590 465738
rect 603970 465418 604002 465654
rect 604238 465418 604322 465654
rect 604558 465418 604590 465654
rect 603970 425974 604590 465418
rect 603970 425738 604002 425974
rect 604238 425738 604322 425974
rect 604558 425738 604590 425974
rect 603970 425654 604590 425738
rect 603970 425418 604002 425654
rect 604238 425418 604322 425654
rect 604558 425418 604590 425654
rect 603970 385974 604590 425418
rect 603970 385738 604002 385974
rect 604238 385738 604322 385974
rect 604558 385738 604590 385974
rect 603970 385654 604590 385738
rect 603970 385418 604002 385654
rect 604238 385418 604322 385654
rect 604558 385418 604590 385654
rect 603970 345974 604590 385418
rect 603970 345738 604002 345974
rect 604238 345738 604322 345974
rect 604558 345738 604590 345974
rect 603970 345654 604590 345738
rect 603970 345418 604002 345654
rect 604238 345418 604322 345654
rect 604558 345418 604590 345654
rect 603970 305974 604590 345418
rect 603970 305738 604002 305974
rect 604238 305738 604322 305974
rect 604558 305738 604590 305974
rect 603970 305654 604590 305738
rect 603970 305418 604002 305654
rect 604238 305418 604322 305654
rect 604558 305418 604590 305654
rect 603970 265974 604590 305418
rect 603970 265738 604002 265974
rect 604238 265738 604322 265974
rect 604558 265738 604590 265974
rect 603970 265654 604590 265738
rect 603970 265418 604002 265654
rect 604238 265418 604322 265654
rect 604558 265418 604590 265654
rect 603970 225974 604590 265418
rect 603970 225738 604002 225974
rect 604238 225738 604322 225974
rect 604558 225738 604590 225974
rect 603970 225654 604590 225738
rect 603970 225418 604002 225654
rect 604238 225418 604322 225654
rect 604558 225418 604590 225654
rect 603970 185974 604590 225418
rect 603970 185738 604002 185974
rect 604238 185738 604322 185974
rect 604558 185738 604590 185974
rect 603970 185654 604590 185738
rect 603970 185418 604002 185654
rect 604238 185418 604322 185654
rect 604558 185418 604590 185654
rect 603970 145974 604590 185418
rect 603970 145738 604002 145974
rect 604238 145738 604322 145974
rect 604558 145738 604590 145974
rect 603970 145654 604590 145738
rect 603970 145418 604002 145654
rect 604238 145418 604322 145654
rect 604558 145418 604590 145654
rect 603970 105974 604590 145418
rect 603970 105738 604002 105974
rect 604238 105738 604322 105974
rect 604558 105738 604590 105974
rect 603970 105654 604590 105738
rect 603970 105418 604002 105654
rect 604238 105418 604322 105654
rect 604558 105418 604590 105654
rect 603970 65974 604590 105418
rect 603970 65738 604002 65974
rect 604238 65738 604322 65974
rect 604558 65738 604590 65974
rect 603970 65654 604590 65738
rect 603970 65418 604002 65654
rect 604238 65418 604322 65654
rect 604558 65418 604590 65654
rect 603970 25974 604590 65418
rect 603970 25738 604002 25974
rect 604238 25738 604322 25974
rect 604558 25738 604590 25974
rect 603970 25654 604590 25738
rect 603970 25418 604002 25654
rect 604238 25418 604322 25654
rect 604558 25418 604590 25654
rect 603970 -19006 604590 25418
rect 603970 -19242 604002 -19006
rect 604238 -19242 604322 -19006
rect 604558 -19242 604590 -19006
rect 603970 -19326 604590 -19242
rect 603970 -19562 604002 -19326
rect 604238 -19562 604322 -19326
rect 604558 -19562 604590 -19326
rect 603970 -19594 604590 -19562
rect 607080 669694 607700 726052
rect 607080 669458 607112 669694
rect 607348 669458 607432 669694
rect 607668 669458 607700 669694
rect 607080 669374 607700 669458
rect 607080 669138 607112 669374
rect 607348 669138 607432 669374
rect 607668 669138 607700 669374
rect 607080 629694 607700 669138
rect 607080 629458 607112 629694
rect 607348 629458 607432 629694
rect 607668 629458 607700 629694
rect 607080 629374 607700 629458
rect 607080 629138 607112 629374
rect 607348 629138 607432 629374
rect 607668 629138 607700 629374
rect 607080 589694 607700 629138
rect 607080 589458 607112 589694
rect 607348 589458 607432 589694
rect 607668 589458 607700 589694
rect 607080 589374 607700 589458
rect 607080 589138 607112 589374
rect 607348 589138 607432 589374
rect 607668 589138 607700 589374
rect 607080 549694 607700 589138
rect 607080 549458 607112 549694
rect 607348 549458 607432 549694
rect 607668 549458 607700 549694
rect 607080 549374 607700 549458
rect 607080 549138 607112 549374
rect 607348 549138 607432 549374
rect 607668 549138 607700 549374
rect 607080 509694 607700 549138
rect 607080 509458 607112 509694
rect 607348 509458 607432 509694
rect 607668 509458 607700 509694
rect 607080 509374 607700 509458
rect 607080 509138 607112 509374
rect 607348 509138 607432 509374
rect 607668 509138 607700 509374
rect 607080 469694 607700 509138
rect 607080 469458 607112 469694
rect 607348 469458 607432 469694
rect 607668 469458 607700 469694
rect 607080 469374 607700 469458
rect 607080 469138 607112 469374
rect 607348 469138 607432 469374
rect 607668 469138 607700 469374
rect 607080 429694 607700 469138
rect 607080 429458 607112 429694
rect 607348 429458 607432 429694
rect 607668 429458 607700 429694
rect 607080 429374 607700 429458
rect 607080 429138 607112 429374
rect 607348 429138 607432 429374
rect 607668 429138 607700 429374
rect 607080 389694 607700 429138
rect 607080 389458 607112 389694
rect 607348 389458 607432 389694
rect 607668 389458 607700 389694
rect 607080 389374 607700 389458
rect 607080 389138 607112 389374
rect 607348 389138 607432 389374
rect 607668 389138 607700 389374
rect 607080 349694 607700 389138
rect 607080 349458 607112 349694
rect 607348 349458 607432 349694
rect 607668 349458 607700 349694
rect 607080 349374 607700 349458
rect 607080 349138 607112 349374
rect 607348 349138 607432 349374
rect 607668 349138 607700 349374
rect 607080 309694 607700 349138
rect 607080 309458 607112 309694
rect 607348 309458 607432 309694
rect 607668 309458 607700 309694
rect 607080 309374 607700 309458
rect 607080 309138 607112 309374
rect 607348 309138 607432 309374
rect 607668 309138 607700 309374
rect 607080 269694 607700 309138
rect 607080 269458 607112 269694
rect 607348 269458 607432 269694
rect 607668 269458 607700 269694
rect 607080 269374 607700 269458
rect 607080 269138 607112 269374
rect 607348 269138 607432 269374
rect 607668 269138 607700 269374
rect 607080 229694 607700 269138
rect 607080 229458 607112 229694
rect 607348 229458 607432 229694
rect 607668 229458 607700 229694
rect 607080 229374 607700 229458
rect 607080 229138 607112 229374
rect 607348 229138 607432 229374
rect 607668 229138 607700 229374
rect 607080 189694 607700 229138
rect 607080 189458 607112 189694
rect 607348 189458 607432 189694
rect 607668 189458 607700 189694
rect 607080 189374 607700 189458
rect 607080 189138 607112 189374
rect 607348 189138 607432 189374
rect 607668 189138 607700 189374
rect 607080 149694 607700 189138
rect 607080 149458 607112 149694
rect 607348 149458 607432 149694
rect 607668 149458 607700 149694
rect 607080 149374 607700 149458
rect 607080 149138 607112 149374
rect 607348 149138 607432 149374
rect 607668 149138 607700 149374
rect 607080 109694 607700 149138
rect 607080 109458 607112 109694
rect 607348 109458 607432 109694
rect 607668 109458 607700 109694
rect 607080 109374 607700 109458
rect 607080 109138 607112 109374
rect 607348 109138 607432 109374
rect 607668 109138 607700 109374
rect 607080 69694 607700 109138
rect 607080 69458 607112 69694
rect 607348 69458 607432 69694
rect 607668 69458 607700 69694
rect 607080 69374 607700 69458
rect 607080 69138 607112 69374
rect 607348 69138 607432 69374
rect 607668 69138 607700 69374
rect 607080 29694 607700 69138
rect 607080 29458 607112 29694
rect 607348 29458 607432 29694
rect 607668 29458 607700 29694
rect 607080 29374 607700 29458
rect 607080 29138 607112 29374
rect 607348 29138 607432 29374
rect 607668 29138 607700 29374
rect 607080 -22116 607700 29138
rect 607080 -22352 607112 -22116
rect 607348 -22352 607432 -22116
rect 607668 -22352 607700 -22116
rect 607080 -22436 607700 -22352
rect 607080 -22672 607112 -22436
rect 607348 -22672 607432 -22436
rect 607668 -22672 607700 -22436
rect 607080 -22704 607700 -22672
<< via4 >>
rect -23744 726372 -23508 726608
rect -23424 726372 -23188 726608
rect -23744 726052 -23508 726288
rect -23424 726052 -23188 726288
rect -23744 669458 -23508 669694
rect -23424 669458 -23188 669694
rect -23744 669138 -23508 669374
rect -23424 669138 -23188 669374
rect -23744 629458 -23508 629694
rect -23424 629458 -23188 629694
rect -23744 629138 -23508 629374
rect -23424 629138 -23188 629374
rect -23744 589458 -23508 589694
rect -23424 589458 -23188 589694
rect -23744 589138 -23508 589374
rect -23424 589138 -23188 589374
rect -23744 549458 -23508 549694
rect -23424 549458 -23188 549694
rect -23744 549138 -23508 549374
rect -23424 549138 -23188 549374
rect -23744 509458 -23508 509694
rect -23424 509458 -23188 509694
rect -23744 509138 -23508 509374
rect -23424 509138 -23188 509374
rect -23744 469458 -23508 469694
rect -23424 469458 -23188 469694
rect -23744 469138 -23508 469374
rect -23424 469138 -23188 469374
rect -23744 429458 -23508 429694
rect -23424 429458 -23188 429694
rect -23744 429138 -23508 429374
rect -23424 429138 -23188 429374
rect -23744 389458 -23508 389694
rect -23424 389458 -23188 389694
rect -23744 389138 -23508 389374
rect -23424 389138 -23188 389374
rect -23744 349458 -23508 349694
rect -23424 349458 -23188 349694
rect -23744 349138 -23508 349374
rect -23424 349138 -23188 349374
rect -23744 309458 -23508 309694
rect -23424 309458 -23188 309694
rect -23744 309138 -23508 309374
rect -23424 309138 -23188 309374
rect -23744 269458 -23508 269694
rect -23424 269458 -23188 269694
rect -23744 269138 -23508 269374
rect -23424 269138 -23188 269374
rect -23744 229458 -23508 229694
rect -23424 229458 -23188 229694
rect -23744 229138 -23508 229374
rect -23424 229138 -23188 229374
rect -23744 189458 -23508 189694
rect -23424 189458 -23188 189694
rect -23744 189138 -23508 189374
rect -23424 189138 -23188 189374
rect -23744 149458 -23508 149694
rect -23424 149458 -23188 149694
rect -23744 149138 -23508 149374
rect -23424 149138 -23188 149374
rect -23744 109458 -23508 109694
rect -23424 109458 -23188 109694
rect -23744 109138 -23508 109374
rect -23424 109138 -23188 109374
rect -23744 69458 -23508 69694
rect -23424 69458 -23188 69694
rect -23744 69138 -23508 69374
rect -23424 69138 -23188 69374
rect -23744 29458 -23508 29694
rect -23424 29458 -23188 29694
rect -23744 29138 -23508 29374
rect -23424 29138 -23188 29374
rect -20634 723262 -20398 723498
rect -20314 723262 -20078 723498
rect -20634 722942 -20398 723178
rect -20314 722942 -20078 723178
rect -20634 665738 -20398 665974
rect -20314 665738 -20078 665974
rect -20634 665418 -20398 665654
rect -20314 665418 -20078 665654
rect -20634 625738 -20398 625974
rect -20314 625738 -20078 625974
rect -20634 625418 -20398 625654
rect -20314 625418 -20078 625654
rect -20634 585738 -20398 585974
rect -20314 585738 -20078 585974
rect -20634 585418 -20398 585654
rect -20314 585418 -20078 585654
rect -20634 545738 -20398 545974
rect -20314 545738 -20078 545974
rect -20634 545418 -20398 545654
rect -20314 545418 -20078 545654
rect -20634 505738 -20398 505974
rect -20314 505738 -20078 505974
rect -20634 505418 -20398 505654
rect -20314 505418 -20078 505654
rect -20634 465738 -20398 465974
rect -20314 465738 -20078 465974
rect -20634 465418 -20398 465654
rect -20314 465418 -20078 465654
rect -20634 425738 -20398 425974
rect -20314 425738 -20078 425974
rect -20634 425418 -20398 425654
rect -20314 425418 -20078 425654
rect -20634 385738 -20398 385974
rect -20314 385738 -20078 385974
rect -20634 385418 -20398 385654
rect -20314 385418 -20078 385654
rect -20634 345738 -20398 345974
rect -20314 345738 -20078 345974
rect -20634 345418 -20398 345654
rect -20314 345418 -20078 345654
rect -20634 305738 -20398 305974
rect -20314 305738 -20078 305974
rect -20634 305418 -20398 305654
rect -20314 305418 -20078 305654
rect -20634 265738 -20398 265974
rect -20314 265738 -20078 265974
rect -20634 265418 -20398 265654
rect -20314 265418 -20078 265654
rect -20634 225738 -20398 225974
rect -20314 225738 -20078 225974
rect -20634 225418 -20398 225654
rect -20314 225418 -20078 225654
rect -20634 185738 -20398 185974
rect -20314 185738 -20078 185974
rect -20634 185418 -20398 185654
rect -20314 185418 -20078 185654
rect -20634 145738 -20398 145974
rect -20314 145738 -20078 145974
rect -20634 145418 -20398 145654
rect -20314 145418 -20078 145654
rect -20634 105738 -20398 105974
rect -20314 105738 -20078 105974
rect -20634 105418 -20398 105654
rect -20314 105418 -20078 105654
rect -20634 65738 -20398 65974
rect -20314 65738 -20078 65974
rect -20634 65418 -20398 65654
rect -20314 65418 -20078 65654
rect -20634 25738 -20398 25974
rect -20314 25738 -20078 25974
rect -20634 25418 -20398 25654
rect -20314 25418 -20078 25654
rect -17524 720152 -17288 720388
rect -17204 720152 -16968 720388
rect -17524 719832 -17288 720068
rect -17204 719832 -16968 720068
rect 607112 726372 607348 726608
rect 607432 726372 607668 726608
rect 607112 726052 607348 726288
rect 607432 726052 607668 726288
rect 604002 723262 604238 723498
rect 604322 723262 604558 723498
rect 604002 722942 604238 723178
rect 604322 722942 604558 723178
rect 580626 720152 580862 720388
rect 580946 720152 581182 720388
rect 580626 719832 580862 720068
rect 580946 719832 581182 720068
rect -17524 662018 -17288 662254
rect -17204 662018 -16968 662254
rect -17524 661698 -17288 661934
rect -17204 661698 -16968 661934
rect -17524 622018 -17288 622254
rect -17204 622018 -16968 622254
rect -17524 621698 -17288 621934
rect -17204 621698 -16968 621934
rect -17524 582018 -17288 582254
rect -17204 582018 -16968 582254
rect -17524 581698 -17288 581934
rect -17204 581698 -16968 581934
rect -17524 542018 -17288 542254
rect -17204 542018 -16968 542254
rect -17524 541698 -17288 541934
rect -17204 541698 -16968 541934
rect -17524 502018 -17288 502254
rect -17204 502018 -16968 502254
rect -17524 501698 -17288 501934
rect -17204 501698 -16968 501934
rect -17524 462018 -17288 462254
rect -17204 462018 -16968 462254
rect -17524 461698 -17288 461934
rect -17204 461698 -16968 461934
rect -17524 422018 -17288 422254
rect -17204 422018 -16968 422254
rect -17524 421698 -17288 421934
rect -17204 421698 -16968 421934
rect -17524 382018 -17288 382254
rect -17204 382018 -16968 382254
rect -17524 381698 -17288 381934
rect -17204 381698 -16968 381934
rect -17524 342018 -17288 342254
rect -17204 342018 -16968 342254
rect -17524 341698 -17288 341934
rect -17204 341698 -16968 341934
rect -17524 302018 -17288 302254
rect -17204 302018 -16968 302254
rect -17524 301698 -17288 301934
rect -17204 301698 -16968 301934
rect -17524 262018 -17288 262254
rect -17204 262018 -16968 262254
rect -17524 261698 -17288 261934
rect -17204 261698 -16968 261934
rect -17524 222018 -17288 222254
rect -17204 222018 -16968 222254
rect -17524 221698 -17288 221934
rect -17204 221698 -16968 221934
rect -17524 182018 -17288 182254
rect -17204 182018 -16968 182254
rect -17524 181698 -17288 181934
rect -17204 181698 -16968 181934
rect -17524 142018 -17288 142254
rect -17204 142018 -16968 142254
rect -17524 141698 -17288 141934
rect -17204 141698 -16968 141934
rect -17524 102018 -17288 102254
rect -17204 102018 -16968 102254
rect -17524 101698 -17288 101934
rect -17204 101698 -16968 101934
rect -17524 62018 -17288 62254
rect -17204 62018 -16968 62254
rect -17524 61698 -17288 61934
rect -17204 61698 -16968 61934
rect -17524 22018 -17288 22254
rect -17204 22018 -16968 22254
rect -17524 21698 -17288 21934
rect -17204 21698 -16968 21934
rect -14414 717042 -14178 717278
rect -14094 717042 -13858 717278
rect -14414 716722 -14178 716958
rect -14094 716722 -13858 716958
rect -14414 698298 -14178 698534
rect -14094 698298 -13858 698534
rect -14414 697978 -14178 698214
rect -14094 697978 -13858 698214
rect -14414 658298 -14178 658534
rect -14094 658298 -13858 658534
rect -14414 657978 -14178 658214
rect -14094 657978 -13858 658214
rect -14414 618298 -14178 618534
rect -14094 618298 -13858 618534
rect -14414 617978 -14178 618214
rect -14094 617978 -13858 618214
rect -14414 578298 -14178 578534
rect -14094 578298 -13858 578534
rect -14414 577978 -14178 578214
rect -14094 577978 -13858 578214
rect -14414 538298 -14178 538534
rect -14094 538298 -13858 538534
rect -14414 537978 -14178 538214
rect -14094 537978 -13858 538214
rect -14414 498298 -14178 498534
rect -14094 498298 -13858 498534
rect -14414 497978 -14178 498214
rect -14094 497978 -13858 498214
rect -14414 458298 -14178 458534
rect -14094 458298 -13858 458534
rect -14414 457978 -14178 458214
rect -14094 457978 -13858 458214
rect -14414 418298 -14178 418534
rect -14094 418298 -13858 418534
rect -14414 417978 -14178 418214
rect -14094 417978 -13858 418214
rect -14414 378298 -14178 378534
rect -14094 378298 -13858 378534
rect -14414 377978 -14178 378214
rect -14094 377978 -13858 378214
rect -14414 338298 -14178 338534
rect -14094 338298 -13858 338534
rect -14414 337978 -14178 338214
rect -14094 337978 -13858 338214
rect -14414 298298 -14178 298534
rect -14094 298298 -13858 298534
rect -14414 297978 -14178 298214
rect -14094 297978 -13858 298214
rect -14414 258298 -14178 258534
rect -14094 258298 -13858 258534
rect -14414 257978 -14178 258214
rect -14094 257978 -13858 258214
rect -14414 218298 -14178 218534
rect -14094 218298 -13858 218534
rect -14414 217978 -14178 218214
rect -14094 217978 -13858 218214
rect -14414 178298 -14178 178534
rect -14094 178298 -13858 178534
rect -14414 177978 -14178 178214
rect -14094 177978 -13858 178214
rect -14414 138298 -14178 138534
rect -14094 138298 -13858 138534
rect -14414 137978 -14178 138214
rect -14094 137978 -13858 138214
rect -14414 98298 -14178 98534
rect -14094 98298 -13858 98534
rect -14414 97978 -14178 98214
rect -14094 97978 -13858 98214
rect -14414 58298 -14178 58534
rect -14094 58298 -13858 58534
rect -14414 57978 -14178 58214
rect -14094 57978 -13858 58214
rect -14414 18298 -14178 18534
rect -14094 18298 -13858 18534
rect -14414 17978 -14178 18214
rect -14094 17978 -13858 18214
rect -11304 713932 -11068 714168
rect -10984 713932 -10748 714168
rect -11304 713612 -11068 713848
rect -10984 713612 -10748 713848
rect -11304 694578 -11068 694814
rect -10984 694578 -10748 694814
rect -11304 694258 -11068 694494
rect -10984 694258 -10748 694494
rect -11304 654578 -11068 654814
rect -10984 654578 -10748 654814
rect -11304 654258 -11068 654494
rect -10984 654258 -10748 654494
rect -11304 614578 -11068 614814
rect -10984 614578 -10748 614814
rect -11304 614258 -11068 614494
rect -10984 614258 -10748 614494
rect -11304 574578 -11068 574814
rect -10984 574578 -10748 574814
rect -11304 574258 -11068 574494
rect -10984 574258 -10748 574494
rect -11304 534578 -11068 534814
rect -10984 534578 -10748 534814
rect -11304 534258 -11068 534494
rect -10984 534258 -10748 534494
rect -11304 494578 -11068 494814
rect -10984 494578 -10748 494814
rect -11304 494258 -11068 494494
rect -10984 494258 -10748 494494
rect -11304 454578 -11068 454814
rect -10984 454578 -10748 454814
rect -11304 454258 -11068 454494
rect -10984 454258 -10748 454494
rect -11304 414578 -11068 414814
rect -10984 414578 -10748 414814
rect -11304 414258 -11068 414494
rect -10984 414258 -10748 414494
rect -11304 374578 -11068 374814
rect -10984 374578 -10748 374814
rect -11304 374258 -11068 374494
rect -10984 374258 -10748 374494
rect -11304 334578 -11068 334814
rect -10984 334578 -10748 334814
rect -11304 334258 -11068 334494
rect -10984 334258 -10748 334494
rect -11304 294578 -11068 294814
rect -10984 294578 -10748 294814
rect -11304 294258 -11068 294494
rect -10984 294258 -10748 294494
rect -11304 254578 -11068 254814
rect -10984 254578 -10748 254814
rect -11304 254258 -11068 254494
rect -10984 254258 -10748 254494
rect -11304 214578 -11068 214814
rect -10984 214578 -10748 214814
rect -11304 214258 -11068 214494
rect -10984 214258 -10748 214494
rect -11304 174578 -11068 174814
rect -10984 174578 -10748 174814
rect -11304 174258 -11068 174494
rect -10984 174258 -10748 174494
rect -11304 134578 -11068 134814
rect -10984 134578 -10748 134814
rect -11304 134258 -11068 134494
rect -10984 134258 -10748 134494
rect -11304 94578 -11068 94814
rect -10984 94578 -10748 94814
rect -11304 94258 -11068 94494
rect -10984 94258 -10748 94494
rect -11304 54578 -11068 54814
rect -10984 54578 -10748 54814
rect -11304 54258 -11068 54494
rect -10984 54258 -10748 54494
rect -11304 14578 -11068 14814
rect -10984 14578 -10748 14814
rect -11304 14258 -11068 14494
rect -10984 14258 -10748 14494
rect -8194 710822 -7958 711058
rect -7874 710822 -7638 711058
rect -8194 710502 -7958 710738
rect -7874 710502 -7638 710738
rect -8194 690858 -7958 691094
rect -7874 690858 -7638 691094
rect -8194 690538 -7958 690774
rect -7874 690538 -7638 690774
rect -8194 650858 -7958 651094
rect -7874 650858 -7638 651094
rect -8194 650538 -7958 650774
rect -7874 650538 -7638 650774
rect -8194 610858 -7958 611094
rect -7874 610858 -7638 611094
rect -8194 610538 -7958 610774
rect -7874 610538 -7638 610774
rect -8194 570858 -7958 571094
rect -7874 570858 -7638 571094
rect -8194 570538 -7958 570774
rect -7874 570538 -7638 570774
rect -8194 530858 -7958 531094
rect -7874 530858 -7638 531094
rect -8194 530538 -7958 530774
rect -7874 530538 -7638 530774
rect -8194 490858 -7958 491094
rect -7874 490858 -7638 491094
rect -8194 490538 -7958 490774
rect -7874 490538 -7638 490774
rect -8194 450858 -7958 451094
rect -7874 450858 -7638 451094
rect -8194 450538 -7958 450774
rect -7874 450538 -7638 450774
rect -8194 410858 -7958 411094
rect -7874 410858 -7638 411094
rect -8194 410538 -7958 410774
rect -7874 410538 -7638 410774
rect -8194 370858 -7958 371094
rect -7874 370858 -7638 371094
rect -8194 370538 -7958 370774
rect -7874 370538 -7638 370774
rect -8194 330858 -7958 331094
rect -7874 330858 -7638 331094
rect -8194 330538 -7958 330774
rect -7874 330538 -7638 330774
rect -8194 290858 -7958 291094
rect -7874 290858 -7638 291094
rect -8194 290538 -7958 290774
rect -7874 290538 -7638 290774
rect -8194 250858 -7958 251094
rect -7874 250858 -7638 251094
rect -8194 250538 -7958 250774
rect -7874 250538 -7638 250774
rect -8194 210858 -7958 211094
rect -7874 210858 -7638 211094
rect -8194 210538 -7958 210774
rect -7874 210538 -7638 210774
rect -8194 170858 -7958 171094
rect -7874 170858 -7638 171094
rect -8194 170538 -7958 170774
rect -7874 170538 -7638 170774
rect -8194 130858 -7958 131094
rect -7874 130858 -7638 131094
rect -8194 130538 -7958 130774
rect -7874 130538 -7638 130774
rect -8194 90858 -7958 91094
rect -7874 90858 -7638 91094
rect -8194 90538 -7958 90774
rect -7874 90538 -7638 90774
rect -8194 50858 -7958 51094
rect -7874 50858 -7638 51094
rect -8194 50538 -7958 50774
rect -7874 50538 -7638 50774
rect -8194 10858 -7958 11094
rect -7874 10858 -7638 11094
rect -8194 10538 -7958 10774
rect -7874 10538 -7638 10774
rect -5084 707712 -4848 707948
rect -4764 707712 -4528 707948
rect -5084 707392 -4848 707628
rect -4764 707392 -4528 707628
rect -5084 687138 -4848 687374
rect -4764 687138 -4528 687374
rect -5084 686818 -4848 687054
rect -4764 686818 -4528 687054
rect -5084 647138 -4848 647374
rect -4764 647138 -4528 647374
rect -5084 646818 -4848 647054
rect -4764 646818 -4528 647054
rect -5084 607138 -4848 607374
rect -4764 607138 -4528 607374
rect -5084 606818 -4848 607054
rect -4764 606818 -4528 607054
rect -5084 567138 -4848 567374
rect -4764 567138 -4528 567374
rect -5084 566818 -4848 567054
rect -4764 566818 -4528 567054
rect -5084 527138 -4848 527374
rect -4764 527138 -4528 527374
rect -5084 526818 -4848 527054
rect -4764 526818 -4528 527054
rect -5084 487138 -4848 487374
rect -4764 487138 -4528 487374
rect -5084 486818 -4848 487054
rect -4764 486818 -4528 487054
rect -5084 447138 -4848 447374
rect -4764 447138 -4528 447374
rect -5084 446818 -4848 447054
rect -4764 446818 -4528 447054
rect -5084 407138 -4848 407374
rect -4764 407138 -4528 407374
rect -5084 406818 -4848 407054
rect -4764 406818 -4528 407054
rect -5084 367138 -4848 367374
rect -4764 367138 -4528 367374
rect -5084 366818 -4848 367054
rect -4764 366818 -4528 367054
rect -5084 327138 -4848 327374
rect -4764 327138 -4528 327374
rect -5084 326818 -4848 327054
rect -4764 326818 -4528 327054
rect -5084 287138 -4848 287374
rect -4764 287138 -4528 287374
rect -5084 286818 -4848 287054
rect -4764 286818 -4528 287054
rect -5084 247138 -4848 247374
rect -4764 247138 -4528 247374
rect -5084 246818 -4848 247054
rect -4764 246818 -4528 247054
rect -5084 207138 -4848 207374
rect -4764 207138 -4528 207374
rect -5084 206818 -4848 207054
rect -4764 206818 -4528 207054
rect -5084 167138 -4848 167374
rect -4764 167138 -4528 167374
rect -5084 166818 -4848 167054
rect -4764 166818 -4528 167054
rect -5084 127138 -4848 127374
rect -4764 127138 -4528 127374
rect -5084 126818 -4848 127054
rect -4764 126818 -4528 127054
rect -5084 87138 -4848 87374
rect -4764 87138 -4528 87374
rect -5084 86818 -4848 87054
rect -4764 86818 -4528 87054
rect -5084 47138 -4848 47374
rect -4764 47138 -4528 47374
rect -5084 46818 -4848 47054
rect -4764 46818 -4528 47054
rect -5084 7138 -4848 7374
rect -4764 7138 -4528 7374
rect -5084 6818 -4848 7054
rect -4764 6818 -4528 7054
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect 7876 693480 8112 693716
rect 8196 693480 8432 693716
rect 7876 693160 8112 693396
rect 8196 693160 8432 693396
rect 38032 693480 38268 693716
rect 38352 693480 38588 693716
rect 38032 693160 38268 693396
rect 38352 693160 38588 693396
rect 74032 693480 74268 693716
rect 74352 693480 74588 693716
rect 74032 693160 74268 693396
rect 74352 693160 74588 693396
rect 110032 693480 110268 693716
rect 110352 693480 110588 693716
rect 110032 693160 110268 693396
rect 110352 693160 110588 693396
rect 146032 693480 146268 693716
rect 146352 693480 146588 693716
rect 146032 693160 146268 693396
rect 146352 693160 146588 693396
rect 182032 693480 182268 693716
rect 182352 693480 182588 693716
rect 182032 693160 182268 693396
rect 182352 693160 182588 693396
rect 218032 693480 218268 693716
rect 218352 693480 218588 693716
rect 218032 693160 218268 693396
rect 218352 693160 218588 693396
rect 254032 693480 254268 693716
rect 254352 693480 254588 693716
rect 254032 693160 254268 693396
rect 254352 693160 254588 693396
rect 290032 693480 290268 693716
rect 290352 693480 290588 693716
rect 290032 693160 290268 693396
rect 290352 693160 290588 693396
rect 326032 693480 326268 693716
rect 326352 693480 326588 693716
rect 326032 693160 326268 693396
rect 326352 693160 326588 693396
rect 362032 693480 362268 693716
rect 362352 693480 362588 693716
rect 362032 693160 362268 693396
rect 362352 693160 362588 693396
rect 398032 693480 398268 693716
rect 398352 693480 398588 693716
rect 398032 693160 398268 693396
rect 398352 693160 398588 693396
rect 434032 693480 434268 693716
rect 434352 693480 434588 693716
rect 434032 693160 434268 693396
rect 434352 693160 434588 693396
rect 470032 693480 470268 693716
rect 470352 693480 470588 693716
rect 470032 693160 470268 693396
rect 470352 693160 470588 693396
rect 506032 693480 506268 693716
rect 506352 693480 506588 693716
rect 506032 693160 506268 693396
rect 506352 693160 506588 693396
rect 542032 693480 542268 693716
rect 542352 693480 542588 693716
rect 542032 693160 542268 693396
rect 542352 693160 542588 693396
rect 571532 693480 571768 693716
rect 571852 693480 572088 693716
rect 571532 693160 571768 693396
rect 571852 693160 572088 693396
rect 9116 692240 9352 692476
rect 9436 692240 9672 692476
rect 9116 691920 9352 692156
rect 9436 691920 9672 692156
rect 56652 692240 56888 692476
rect 56972 692240 57208 692476
rect 56652 691920 56888 692156
rect 56972 691920 57208 692156
rect 92652 692240 92888 692476
rect 92972 692240 93208 692476
rect 92652 691920 92888 692156
rect 92972 691920 93208 692156
rect 128652 692240 128888 692476
rect 128972 692240 129208 692476
rect 128652 691920 128888 692156
rect 128972 691920 129208 692156
rect 164652 692240 164888 692476
rect 164972 692240 165208 692476
rect 164652 691920 164888 692156
rect 164972 691920 165208 692156
rect 200652 692240 200888 692476
rect 200972 692240 201208 692476
rect 200652 691920 200888 692156
rect 200972 691920 201208 692156
rect 236652 692240 236888 692476
rect 236972 692240 237208 692476
rect 236652 691920 236888 692156
rect 236972 691920 237208 692156
rect 272652 692240 272888 692476
rect 272972 692240 273208 692476
rect 272652 691920 272888 692156
rect 272972 691920 273208 692156
rect 308652 692240 308888 692476
rect 308972 692240 309208 692476
rect 308652 691920 308888 692156
rect 308972 691920 309208 692156
rect 344652 692240 344888 692476
rect 344972 692240 345208 692476
rect 344652 691920 344888 692156
rect 344972 691920 345208 692156
rect 380652 692240 380888 692476
rect 380972 692240 381208 692476
rect 380652 691920 380888 692156
rect 380972 691920 381208 692156
rect 416652 692240 416888 692476
rect 416972 692240 417208 692476
rect 416652 691920 416888 692156
rect 416972 691920 417208 692156
rect 452652 692240 452888 692476
rect 452972 692240 453208 692476
rect 452652 691920 452888 692156
rect 452972 691920 453208 692156
rect 488652 692240 488888 692476
rect 488972 692240 489208 692476
rect 488652 691920 488888 692156
rect 488972 691920 489208 692156
rect 524652 692240 524888 692476
rect 524972 692240 525208 692476
rect 524652 691920 524888 692156
rect 524972 691920 525208 692156
rect 560652 692240 560888 692476
rect 560972 692240 561208 692476
rect 560652 691920 560888 692156
rect 560972 691920 561208 692156
rect 570292 692240 570528 692476
rect 570612 692240 570848 692476
rect 570292 691920 570528 692156
rect 570612 691920 570848 692156
rect 7876 687138 8112 687374
rect 8196 687138 8432 687374
rect 7876 686818 8112 687054
rect 8196 686818 8432 687054
rect 38032 687138 38268 687374
rect 38352 687138 38588 687374
rect 38032 686818 38268 687054
rect 38352 686818 38588 687054
rect 74032 687138 74268 687374
rect 74352 687138 74588 687374
rect 74032 686818 74268 687054
rect 74352 686818 74588 687054
rect 110032 687138 110268 687374
rect 110352 687138 110588 687374
rect 110032 686818 110268 687054
rect 110352 686818 110588 687054
rect 146032 687138 146268 687374
rect 146352 687138 146588 687374
rect 146032 686818 146268 687054
rect 146352 686818 146588 687054
rect 182032 687138 182268 687374
rect 182352 687138 182588 687374
rect 182032 686818 182268 687054
rect 182352 686818 182588 687054
rect 218032 687138 218268 687374
rect 218352 687138 218588 687374
rect 218032 686818 218268 687054
rect 218352 686818 218588 687054
rect 254032 687138 254268 687374
rect 254352 687138 254588 687374
rect 254032 686818 254268 687054
rect 254352 686818 254588 687054
rect 290032 687138 290268 687374
rect 290352 687138 290588 687374
rect 290032 686818 290268 687054
rect 290352 686818 290588 687054
rect 326032 687138 326268 687374
rect 326352 687138 326588 687374
rect 326032 686818 326268 687054
rect 326352 686818 326588 687054
rect 362032 687138 362268 687374
rect 362352 687138 362588 687374
rect 362032 686818 362268 687054
rect 362352 686818 362588 687054
rect 398032 687138 398268 687374
rect 398352 687138 398588 687374
rect 398032 686818 398268 687054
rect 398352 686818 398588 687054
rect 434032 687138 434268 687374
rect 434352 687138 434588 687374
rect 434032 686818 434268 687054
rect 434352 686818 434588 687054
rect 470032 687138 470268 687374
rect 470352 687138 470588 687374
rect 470032 686818 470268 687054
rect 470352 686818 470588 687054
rect 506032 687138 506268 687374
rect 506352 687138 506588 687374
rect 506032 686818 506268 687054
rect 506352 686818 506588 687054
rect 542032 687138 542268 687374
rect 542352 687138 542588 687374
rect 542032 686818 542268 687054
rect 542352 686818 542588 687054
rect 571532 687138 571768 687374
rect 571852 687138 572088 687374
rect 571532 686818 571768 687054
rect 571852 686818 572088 687054
rect -1974 683418 -1738 683654
rect -1654 683418 -1418 683654
rect -1974 683098 -1738 683334
rect -1654 683098 -1418 683334
rect 9116 683418 9352 683654
rect 9436 683418 9672 683654
rect 9116 683098 9352 683334
rect 9436 683098 9672 683334
rect 56652 683418 56888 683654
rect 56972 683418 57208 683654
rect 56652 683098 56888 683334
rect 56972 683098 57208 683334
rect 92652 683418 92888 683654
rect 92972 683418 93208 683654
rect 92652 683098 92888 683334
rect 92972 683098 93208 683334
rect 128652 683418 128888 683654
rect 128972 683418 129208 683654
rect 128652 683098 128888 683334
rect 128972 683098 129208 683334
rect 164652 683418 164888 683654
rect 164972 683418 165208 683654
rect 164652 683098 164888 683334
rect 164972 683098 165208 683334
rect 200652 683418 200888 683654
rect 200972 683418 201208 683654
rect 200652 683098 200888 683334
rect 200972 683098 201208 683334
rect 236652 683418 236888 683654
rect 236972 683418 237208 683654
rect 236652 683098 236888 683334
rect 236972 683098 237208 683334
rect 272652 683418 272888 683654
rect 272972 683418 273208 683654
rect 272652 683098 272888 683334
rect 272972 683098 273208 683334
rect 308652 683418 308888 683654
rect 308972 683418 309208 683654
rect 308652 683098 308888 683334
rect 308972 683098 309208 683334
rect 344652 683418 344888 683654
rect 344972 683418 345208 683654
rect 344652 683098 344888 683334
rect 344972 683098 345208 683334
rect 380652 683418 380888 683654
rect 380972 683418 381208 683654
rect 380652 683098 380888 683334
rect 380972 683098 381208 683334
rect 416652 683418 416888 683654
rect 416972 683418 417208 683654
rect 416652 683098 416888 683334
rect 416972 683098 417208 683334
rect 452652 683418 452888 683654
rect 452972 683418 453208 683654
rect 452652 683098 452888 683334
rect 452972 683098 453208 683334
rect 488652 683418 488888 683654
rect 488972 683418 489208 683654
rect 488652 683098 488888 683334
rect 488972 683098 489208 683334
rect 524652 683418 524888 683654
rect 524972 683418 525208 683654
rect 524652 683098 524888 683334
rect 524972 683098 525208 683334
rect 560652 683418 560888 683654
rect 560972 683418 561208 683654
rect 560652 683098 560888 683334
rect 560972 683098 561208 683334
rect 570292 683418 570528 683654
rect 570612 683418 570848 683654
rect 570292 683098 570528 683334
rect 570612 683098 570848 683334
rect 600892 720152 601128 720388
rect 601212 720152 601448 720388
rect 600892 719832 601128 720068
rect 601212 719832 601448 720068
rect 597782 717042 598018 717278
rect 598102 717042 598338 717278
rect 597782 716722 598018 716958
rect 598102 716722 598338 716958
rect 594672 713932 594908 714168
rect 594992 713932 595228 714168
rect 594672 713612 594908 713848
rect 594992 713612 595228 713848
rect 591562 710822 591798 711058
rect 591882 710822 592118 711058
rect 591562 710502 591798 710738
rect 591882 710502 592118 710738
rect 588452 707712 588688 707948
rect 588772 707712 589008 707948
rect 588452 707392 588688 707628
rect 588772 707392 589008 707628
rect 580626 662018 580862 662254
rect 580946 662018 581182 662254
rect 580626 661698 580862 661934
rect 580946 661698 581182 661934
rect 7876 647138 8112 647374
rect 8196 647138 8432 647374
rect 7876 646818 8112 647054
rect 8196 646818 8432 647054
rect 38032 647138 38268 647374
rect 38352 647138 38588 647374
rect 38032 646818 38268 647054
rect 38352 646818 38588 647054
rect 74032 647138 74268 647374
rect 74352 647138 74588 647374
rect 74032 646818 74268 647054
rect 74352 646818 74588 647054
rect 110032 647138 110268 647374
rect 110352 647138 110588 647374
rect 110032 646818 110268 647054
rect 110352 646818 110588 647054
rect 146032 647138 146268 647374
rect 146352 647138 146588 647374
rect 146032 646818 146268 647054
rect 146352 646818 146588 647054
rect 182032 647138 182268 647374
rect 182352 647138 182588 647374
rect 182032 646818 182268 647054
rect 182352 646818 182588 647054
rect 218032 647138 218268 647374
rect 218352 647138 218588 647374
rect 218032 646818 218268 647054
rect 218352 646818 218588 647054
rect 254032 647138 254268 647374
rect 254352 647138 254588 647374
rect 254032 646818 254268 647054
rect 254352 646818 254588 647054
rect 290032 647138 290268 647374
rect 290352 647138 290588 647374
rect 290032 646818 290268 647054
rect 290352 646818 290588 647054
rect 326032 647138 326268 647374
rect 326352 647138 326588 647374
rect 326032 646818 326268 647054
rect 326352 646818 326588 647054
rect 362032 647138 362268 647374
rect 362352 647138 362588 647374
rect 362032 646818 362268 647054
rect 362352 646818 362588 647054
rect 398032 647138 398268 647374
rect 398352 647138 398588 647374
rect 398032 646818 398268 647054
rect 398352 646818 398588 647054
rect 434032 647138 434268 647374
rect 434352 647138 434588 647374
rect 434032 646818 434268 647054
rect 434352 646818 434588 647054
rect 470032 647138 470268 647374
rect 470352 647138 470588 647374
rect 470032 646818 470268 647054
rect 470352 646818 470588 647054
rect 506032 647138 506268 647374
rect 506352 647138 506588 647374
rect 506032 646818 506268 647054
rect 506352 646818 506588 647054
rect 542032 647138 542268 647374
rect 542352 647138 542588 647374
rect 542032 646818 542268 647054
rect 542352 646818 542588 647054
rect 571532 647138 571768 647374
rect 571852 647138 572088 647374
rect 571532 646818 571768 647054
rect 571852 646818 572088 647054
rect -1974 643418 -1738 643654
rect -1654 643418 -1418 643654
rect -1974 643098 -1738 643334
rect -1654 643098 -1418 643334
rect 9116 643418 9352 643654
rect 9436 643418 9672 643654
rect 9116 643098 9352 643334
rect 9436 643098 9672 643334
rect 56652 643418 56888 643654
rect 56972 643418 57208 643654
rect 56652 643098 56888 643334
rect 56972 643098 57208 643334
rect 92652 643418 92888 643654
rect 92972 643418 93208 643654
rect 92652 643098 92888 643334
rect 92972 643098 93208 643334
rect 128652 643418 128888 643654
rect 128972 643418 129208 643654
rect 128652 643098 128888 643334
rect 128972 643098 129208 643334
rect 164652 643418 164888 643654
rect 164972 643418 165208 643654
rect 164652 643098 164888 643334
rect 164972 643098 165208 643334
rect 200652 643418 200888 643654
rect 200972 643418 201208 643654
rect 200652 643098 200888 643334
rect 200972 643098 201208 643334
rect 236652 643418 236888 643654
rect 236972 643418 237208 643654
rect 236652 643098 236888 643334
rect 236972 643098 237208 643334
rect 272652 643418 272888 643654
rect 272972 643418 273208 643654
rect 272652 643098 272888 643334
rect 272972 643098 273208 643334
rect 308652 643418 308888 643654
rect 308972 643418 309208 643654
rect 308652 643098 308888 643334
rect 308972 643098 309208 643334
rect 344652 643418 344888 643654
rect 344972 643418 345208 643654
rect 344652 643098 344888 643334
rect 344972 643098 345208 643334
rect 380652 643418 380888 643654
rect 380972 643418 381208 643654
rect 380652 643098 380888 643334
rect 380972 643098 381208 643334
rect 416652 643418 416888 643654
rect 416972 643418 417208 643654
rect 416652 643098 416888 643334
rect 416972 643098 417208 643334
rect 452652 643418 452888 643654
rect 452972 643418 453208 643654
rect 452652 643098 452888 643334
rect 452972 643098 453208 643334
rect 488652 643418 488888 643654
rect 488972 643418 489208 643654
rect 488652 643098 488888 643334
rect 488972 643098 489208 643334
rect 524652 643418 524888 643654
rect 524972 643418 525208 643654
rect 524652 643098 524888 643334
rect 524972 643098 525208 643334
rect 560652 643418 560888 643654
rect 560972 643418 561208 643654
rect 560652 643098 560888 643334
rect 560972 643098 561208 643334
rect 570292 643418 570528 643654
rect 570612 643418 570848 643654
rect 570292 643098 570528 643334
rect 570612 643098 570848 643334
rect 580626 622018 580862 622254
rect 580946 622018 581182 622254
rect 580626 621698 580862 621934
rect 580946 621698 581182 621934
rect 7876 607138 8112 607374
rect 8196 607138 8432 607374
rect 7876 606818 8112 607054
rect 8196 606818 8432 607054
rect 38032 607138 38268 607374
rect 38352 607138 38588 607374
rect 38032 606818 38268 607054
rect 38352 606818 38588 607054
rect 74032 607138 74268 607374
rect 74352 607138 74588 607374
rect 74032 606818 74268 607054
rect 74352 606818 74588 607054
rect 110032 607138 110268 607374
rect 110352 607138 110588 607374
rect 110032 606818 110268 607054
rect 110352 606818 110588 607054
rect 146032 607138 146268 607374
rect 146352 607138 146588 607374
rect 146032 606818 146268 607054
rect 146352 606818 146588 607054
rect 182032 607138 182268 607374
rect 182352 607138 182588 607374
rect 182032 606818 182268 607054
rect 182352 606818 182588 607054
rect 218032 607138 218268 607374
rect 218352 607138 218588 607374
rect 218032 606818 218268 607054
rect 218352 606818 218588 607054
rect 254032 607138 254268 607374
rect 254352 607138 254588 607374
rect 254032 606818 254268 607054
rect 254352 606818 254588 607054
rect 290032 607138 290268 607374
rect 290352 607138 290588 607374
rect 290032 606818 290268 607054
rect 290352 606818 290588 607054
rect 326032 607138 326268 607374
rect 326352 607138 326588 607374
rect 326032 606818 326268 607054
rect 326352 606818 326588 607054
rect 362032 607138 362268 607374
rect 362352 607138 362588 607374
rect 362032 606818 362268 607054
rect 362352 606818 362588 607054
rect 398032 607138 398268 607374
rect 398352 607138 398588 607374
rect 398032 606818 398268 607054
rect 398352 606818 398588 607054
rect 434032 607138 434268 607374
rect 434352 607138 434588 607374
rect 434032 606818 434268 607054
rect 434352 606818 434588 607054
rect 470032 607138 470268 607374
rect 470352 607138 470588 607374
rect 470032 606818 470268 607054
rect 470352 606818 470588 607054
rect 506032 607138 506268 607374
rect 506352 607138 506588 607374
rect 506032 606818 506268 607054
rect 506352 606818 506588 607054
rect 542032 607138 542268 607374
rect 542352 607138 542588 607374
rect 542032 606818 542268 607054
rect 542352 606818 542588 607054
rect 571532 607138 571768 607374
rect 571852 607138 572088 607374
rect 571532 606818 571768 607054
rect 571852 606818 572088 607054
rect -1974 603418 -1738 603654
rect -1654 603418 -1418 603654
rect -1974 603098 -1738 603334
rect -1654 603098 -1418 603334
rect 9116 603418 9352 603654
rect 9436 603418 9672 603654
rect 9116 603098 9352 603334
rect 9436 603098 9672 603334
rect 56652 603418 56888 603654
rect 56972 603418 57208 603654
rect 56652 603098 56888 603334
rect 56972 603098 57208 603334
rect 92652 603418 92888 603654
rect 92972 603418 93208 603654
rect 92652 603098 92888 603334
rect 92972 603098 93208 603334
rect 128652 603418 128888 603654
rect 128972 603418 129208 603654
rect 128652 603098 128888 603334
rect 128972 603098 129208 603334
rect 164652 603418 164888 603654
rect 164972 603418 165208 603654
rect 164652 603098 164888 603334
rect 164972 603098 165208 603334
rect 200652 603418 200888 603654
rect 200972 603418 201208 603654
rect 200652 603098 200888 603334
rect 200972 603098 201208 603334
rect 236652 603418 236888 603654
rect 236972 603418 237208 603654
rect 236652 603098 236888 603334
rect 236972 603098 237208 603334
rect 272652 603418 272888 603654
rect 272972 603418 273208 603654
rect 272652 603098 272888 603334
rect 272972 603098 273208 603334
rect 308652 603418 308888 603654
rect 308972 603418 309208 603654
rect 308652 603098 308888 603334
rect 308972 603098 309208 603334
rect 344652 603418 344888 603654
rect 344972 603418 345208 603654
rect 344652 603098 344888 603334
rect 344972 603098 345208 603334
rect 380652 603418 380888 603654
rect 380972 603418 381208 603654
rect 380652 603098 380888 603334
rect 380972 603098 381208 603334
rect 416652 603418 416888 603654
rect 416972 603418 417208 603654
rect 416652 603098 416888 603334
rect 416972 603098 417208 603334
rect 452652 603418 452888 603654
rect 452972 603418 453208 603654
rect 452652 603098 452888 603334
rect 452972 603098 453208 603334
rect 488652 603418 488888 603654
rect 488972 603418 489208 603654
rect 488652 603098 488888 603334
rect 488972 603098 489208 603334
rect 524652 603418 524888 603654
rect 524972 603418 525208 603654
rect 524652 603098 524888 603334
rect 524972 603098 525208 603334
rect 560652 603418 560888 603654
rect 560972 603418 561208 603654
rect 560652 603098 560888 603334
rect 560972 603098 561208 603334
rect 570292 603418 570528 603654
rect 570612 603418 570848 603654
rect 570292 603098 570528 603334
rect 570612 603098 570848 603334
rect 580626 582018 580862 582254
rect 580946 582018 581182 582254
rect 580626 581698 580862 581934
rect 580946 581698 581182 581934
rect 7876 567138 8112 567374
rect 8196 567138 8432 567374
rect 7876 566818 8112 567054
rect 8196 566818 8432 567054
rect 38032 567138 38268 567374
rect 38352 567138 38588 567374
rect 38032 566818 38268 567054
rect 38352 566818 38588 567054
rect 74032 567138 74268 567374
rect 74352 567138 74588 567374
rect 74032 566818 74268 567054
rect 74352 566818 74588 567054
rect 110032 567138 110268 567374
rect 110352 567138 110588 567374
rect 110032 566818 110268 567054
rect 110352 566818 110588 567054
rect 146032 567138 146268 567374
rect 146352 567138 146588 567374
rect 146032 566818 146268 567054
rect 146352 566818 146588 567054
rect 182032 567138 182268 567374
rect 182352 567138 182588 567374
rect 182032 566818 182268 567054
rect 182352 566818 182588 567054
rect 218032 567138 218268 567374
rect 218352 567138 218588 567374
rect 218032 566818 218268 567054
rect 218352 566818 218588 567054
rect 254032 567138 254268 567374
rect 254352 567138 254588 567374
rect 254032 566818 254268 567054
rect 254352 566818 254588 567054
rect 290032 567138 290268 567374
rect 290352 567138 290588 567374
rect 290032 566818 290268 567054
rect 290352 566818 290588 567054
rect 326032 567138 326268 567374
rect 326352 567138 326588 567374
rect 326032 566818 326268 567054
rect 326352 566818 326588 567054
rect 362032 567138 362268 567374
rect 362352 567138 362588 567374
rect 362032 566818 362268 567054
rect 362352 566818 362588 567054
rect 398032 567138 398268 567374
rect 398352 567138 398588 567374
rect 398032 566818 398268 567054
rect 398352 566818 398588 567054
rect 434032 567138 434268 567374
rect 434352 567138 434588 567374
rect 434032 566818 434268 567054
rect 434352 566818 434588 567054
rect 470032 567138 470268 567374
rect 470352 567138 470588 567374
rect 470032 566818 470268 567054
rect 470352 566818 470588 567054
rect 506032 567138 506268 567374
rect 506352 567138 506588 567374
rect 506032 566818 506268 567054
rect 506352 566818 506588 567054
rect 542032 567138 542268 567374
rect 542352 567138 542588 567374
rect 542032 566818 542268 567054
rect 542352 566818 542588 567054
rect 571532 567138 571768 567374
rect 571852 567138 572088 567374
rect 571532 566818 571768 567054
rect 571852 566818 572088 567054
rect -1974 563418 -1738 563654
rect -1654 563418 -1418 563654
rect -1974 563098 -1738 563334
rect -1654 563098 -1418 563334
rect 9116 563418 9352 563654
rect 9436 563418 9672 563654
rect 9116 563098 9352 563334
rect 9436 563098 9672 563334
rect 56652 563418 56888 563654
rect 56972 563418 57208 563654
rect 56652 563098 56888 563334
rect 56972 563098 57208 563334
rect 92652 563418 92888 563654
rect 92972 563418 93208 563654
rect 92652 563098 92888 563334
rect 92972 563098 93208 563334
rect 128652 563418 128888 563654
rect 128972 563418 129208 563654
rect 128652 563098 128888 563334
rect 128972 563098 129208 563334
rect 164652 563418 164888 563654
rect 164972 563418 165208 563654
rect 164652 563098 164888 563334
rect 164972 563098 165208 563334
rect 200652 563418 200888 563654
rect 200972 563418 201208 563654
rect 200652 563098 200888 563334
rect 200972 563098 201208 563334
rect 236652 563418 236888 563654
rect 236972 563418 237208 563654
rect 236652 563098 236888 563334
rect 236972 563098 237208 563334
rect 272652 563418 272888 563654
rect 272972 563418 273208 563654
rect 272652 563098 272888 563334
rect 272972 563098 273208 563334
rect 308652 563418 308888 563654
rect 308972 563418 309208 563654
rect 308652 563098 308888 563334
rect 308972 563098 309208 563334
rect 344652 563418 344888 563654
rect 344972 563418 345208 563654
rect 344652 563098 344888 563334
rect 344972 563098 345208 563334
rect 380652 563418 380888 563654
rect 380972 563418 381208 563654
rect 380652 563098 380888 563334
rect 380972 563098 381208 563334
rect 416652 563418 416888 563654
rect 416972 563418 417208 563654
rect 416652 563098 416888 563334
rect 416972 563098 417208 563334
rect 452652 563418 452888 563654
rect 452972 563418 453208 563654
rect 452652 563098 452888 563334
rect 452972 563098 453208 563334
rect 488652 563418 488888 563654
rect 488972 563418 489208 563654
rect 488652 563098 488888 563334
rect 488972 563098 489208 563334
rect 524652 563418 524888 563654
rect 524972 563418 525208 563654
rect 524652 563098 524888 563334
rect 524972 563098 525208 563334
rect 560652 563418 560888 563654
rect 560972 563418 561208 563654
rect 560652 563098 560888 563334
rect 560972 563098 561208 563334
rect 570292 563418 570528 563654
rect 570612 563418 570848 563654
rect 570292 563098 570528 563334
rect 570612 563098 570848 563334
rect 580626 542018 580862 542254
rect 580946 542018 581182 542254
rect 580626 541698 580862 541934
rect 580946 541698 581182 541934
rect 7876 527138 8112 527374
rect 8196 527138 8432 527374
rect 7876 526818 8112 527054
rect 8196 526818 8432 527054
rect 38032 527138 38268 527374
rect 38352 527138 38588 527374
rect 38032 526818 38268 527054
rect 38352 526818 38588 527054
rect 74032 527138 74268 527374
rect 74352 527138 74588 527374
rect 74032 526818 74268 527054
rect 74352 526818 74588 527054
rect 110032 527138 110268 527374
rect 110352 527138 110588 527374
rect 110032 526818 110268 527054
rect 110352 526818 110588 527054
rect 146032 527138 146268 527374
rect 146352 527138 146588 527374
rect 146032 526818 146268 527054
rect 146352 526818 146588 527054
rect 182032 527138 182268 527374
rect 182352 527138 182588 527374
rect 182032 526818 182268 527054
rect 182352 526818 182588 527054
rect 218032 527138 218268 527374
rect 218352 527138 218588 527374
rect 218032 526818 218268 527054
rect 218352 526818 218588 527054
rect 254032 527138 254268 527374
rect 254352 527138 254588 527374
rect 254032 526818 254268 527054
rect 254352 526818 254588 527054
rect 290032 527138 290268 527374
rect 290352 527138 290588 527374
rect 290032 526818 290268 527054
rect 290352 526818 290588 527054
rect 326032 527138 326268 527374
rect 326352 527138 326588 527374
rect 326032 526818 326268 527054
rect 326352 526818 326588 527054
rect 362032 527138 362268 527374
rect 362352 527138 362588 527374
rect 362032 526818 362268 527054
rect 362352 526818 362588 527054
rect 398032 527138 398268 527374
rect 398352 527138 398588 527374
rect 398032 526818 398268 527054
rect 398352 526818 398588 527054
rect 434032 527138 434268 527374
rect 434352 527138 434588 527374
rect 434032 526818 434268 527054
rect 434352 526818 434588 527054
rect 470032 527138 470268 527374
rect 470352 527138 470588 527374
rect 470032 526818 470268 527054
rect 470352 526818 470588 527054
rect 506032 527138 506268 527374
rect 506352 527138 506588 527374
rect 506032 526818 506268 527054
rect 506352 526818 506588 527054
rect 542032 527138 542268 527374
rect 542352 527138 542588 527374
rect 542032 526818 542268 527054
rect 542352 526818 542588 527054
rect 571532 527138 571768 527374
rect 571852 527138 572088 527374
rect 571532 526818 571768 527054
rect 571852 526818 572088 527054
rect -1974 523418 -1738 523654
rect -1654 523418 -1418 523654
rect -1974 523098 -1738 523334
rect -1654 523098 -1418 523334
rect 9116 523418 9352 523654
rect 9436 523418 9672 523654
rect 9116 523098 9352 523334
rect 9436 523098 9672 523334
rect 56652 523418 56888 523654
rect 56972 523418 57208 523654
rect 56652 523098 56888 523334
rect 56972 523098 57208 523334
rect 92652 523418 92888 523654
rect 92972 523418 93208 523654
rect 92652 523098 92888 523334
rect 92972 523098 93208 523334
rect 128652 523418 128888 523654
rect 128972 523418 129208 523654
rect 128652 523098 128888 523334
rect 128972 523098 129208 523334
rect 164652 523418 164888 523654
rect 164972 523418 165208 523654
rect 164652 523098 164888 523334
rect 164972 523098 165208 523334
rect 200652 523418 200888 523654
rect 200972 523418 201208 523654
rect 200652 523098 200888 523334
rect 200972 523098 201208 523334
rect 236652 523418 236888 523654
rect 236972 523418 237208 523654
rect 236652 523098 236888 523334
rect 236972 523098 237208 523334
rect 272652 523418 272888 523654
rect 272972 523418 273208 523654
rect 272652 523098 272888 523334
rect 272972 523098 273208 523334
rect 308652 523418 308888 523654
rect 308972 523418 309208 523654
rect 308652 523098 308888 523334
rect 308972 523098 309208 523334
rect 344652 523418 344888 523654
rect 344972 523418 345208 523654
rect 344652 523098 344888 523334
rect 344972 523098 345208 523334
rect 380652 523418 380888 523654
rect 380972 523418 381208 523654
rect 380652 523098 380888 523334
rect 380972 523098 381208 523334
rect 416652 523418 416888 523654
rect 416972 523418 417208 523654
rect 416652 523098 416888 523334
rect 416972 523098 417208 523334
rect 452652 523418 452888 523654
rect 452972 523418 453208 523654
rect 452652 523098 452888 523334
rect 452972 523098 453208 523334
rect 488652 523418 488888 523654
rect 488972 523418 489208 523654
rect 488652 523098 488888 523334
rect 488972 523098 489208 523334
rect 524652 523418 524888 523654
rect 524972 523418 525208 523654
rect 524652 523098 524888 523334
rect 524972 523098 525208 523334
rect 560652 523418 560888 523654
rect 560972 523418 561208 523654
rect 560652 523098 560888 523334
rect 560972 523098 561208 523334
rect 570292 523418 570528 523654
rect 570612 523418 570848 523654
rect 570292 523098 570528 523334
rect 570612 523098 570848 523334
rect 580626 502018 580862 502254
rect 580946 502018 581182 502254
rect 580626 501698 580862 501934
rect 580946 501698 581182 501934
rect 7876 487138 8112 487374
rect 8196 487138 8432 487374
rect 7876 486818 8112 487054
rect 8196 486818 8432 487054
rect 38032 487138 38268 487374
rect 38352 487138 38588 487374
rect 38032 486818 38268 487054
rect 38352 486818 38588 487054
rect 60622 487138 60858 487374
rect 60622 486818 60858 487054
rect 159098 487138 159334 487374
rect 159098 486818 159334 487054
rect 182032 487138 182268 487374
rect 182352 487138 182588 487374
rect 182032 486818 182268 487054
rect 182352 486818 182588 487054
rect 185622 487138 185858 487374
rect 185622 486818 185858 487054
rect 284098 487138 284334 487374
rect 284098 486818 284334 487054
rect 290032 487138 290268 487374
rect 290352 487138 290588 487374
rect 290032 486818 290268 487054
rect 290352 486818 290588 487054
rect 310622 487138 310858 487374
rect 310622 486818 310858 487054
rect 409098 487138 409334 487374
rect 409098 486818 409334 487054
rect 434032 487138 434268 487374
rect 434352 487138 434588 487374
rect 434032 486818 434268 487054
rect 434352 486818 434588 487054
rect 436622 487138 436858 487374
rect 436622 486818 436858 487054
rect 535098 487138 535334 487374
rect 535098 486818 535334 487054
rect 542032 487138 542268 487374
rect 542352 487138 542588 487374
rect 542032 486818 542268 487054
rect 542352 486818 542588 487054
rect 571532 487138 571768 487374
rect 571852 487138 572088 487374
rect 571532 486818 571768 487054
rect 571852 486818 572088 487054
rect -1974 483418 -1738 483654
rect -1654 483418 -1418 483654
rect -1974 483098 -1738 483334
rect -1654 483098 -1418 483334
rect 9116 483418 9352 483654
rect 9436 483418 9672 483654
rect 9116 483098 9352 483334
rect 9436 483098 9672 483334
rect 56652 483418 56888 483654
rect 56972 483418 57208 483654
rect 56652 483098 56888 483334
rect 56972 483098 57208 483334
rect 61342 483418 61578 483654
rect 61342 483098 61578 483334
rect 158378 483418 158614 483654
rect 158378 483098 158614 483334
rect 164652 483418 164888 483654
rect 164972 483418 165208 483654
rect 164652 483098 164888 483334
rect 164972 483098 165208 483334
rect 186342 483418 186578 483654
rect 186342 483098 186578 483334
rect 283378 483418 283614 483654
rect 283378 483098 283614 483334
rect 308652 483418 308888 483654
rect 308972 483418 309208 483654
rect 308652 483098 308888 483334
rect 308972 483098 309208 483334
rect 311342 483418 311578 483654
rect 311342 483098 311578 483334
rect 408378 483418 408614 483654
rect 408378 483098 408614 483334
rect 416652 483418 416888 483654
rect 416972 483418 417208 483654
rect 416652 483098 416888 483334
rect 416972 483098 417208 483334
rect 437342 483418 437578 483654
rect 437342 483098 437578 483334
rect 534378 483418 534614 483654
rect 534378 483098 534614 483334
rect 560652 483418 560888 483654
rect 560972 483418 561208 483654
rect 560652 483098 560888 483334
rect 560972 483098 561208 483334
rect 570292 483418 570528 483654
rect 570612 483418 570848 483654
rect 570292 483098 570528 483334
rect 570612 483098 570848 483334
rect 580626 462018 580862 462254
rect 580946 462018 581182 462254
rect 580626 461698 580862 461934
rect 580946 461698 581182 461934
rect 7876 447138 8112 447374
rect 8196 447138 8432 447374
rect 7876 446818 8112 447054
rect 8196 446818 8432 447054
rect 38032 447138 38268 447374
rect 38352 447138 38588 447374
rect 38032 446818 38268 447054
rect 38352 446818 38588 447054
rect 60622 447138 60858 447374
rect 60622 446818 60858 447054
rect 159098 447138 159334 447374
rect 159098 446818 159334 447054
rect 182032 447138 182268 447374
rect 182352 447138 182588 447374
rect 182032 446818 182268 447054
rect 182352 446818 182588 447054
rect 185622 447138 185858 447374
rect 185622 446818 185858 447054
rect 284098 447138 284334 447374
rect 284098 446818 284334 447054
rect 290032 447138 290268 447374
rect 290352 447138 290588 447374
rect 290032 446818 290268 447054
rect 290352 446818 290588 447054
rect 310622 447138 310858 447374
rect 310622 446818 310858 447054
rect 409098 447138 409334 447374
rect 409098 446818 409334 447054
rect 434032 447138 434268 447374
rect 434352 447138 434588 447374
rect 434032 446818 434268 447054
rect 434352 446818 434588 447054
rect 436622 447138 436858 447374
rect 436622 446818 436858 447054
rect 535098 447138 535334 447374
rect 535098 446818 535334 447054
rect 542032 447138 542268 447374
rect 542352 447138 542588 447374
rect 542032 446818 542268 447054
rect 542352 446818 542588 447054
rect 571532 447138 571768 447374
rect 571852 447138 572088 447374
rect 571532 446818 571768 447054
rect 571852 446818 572088 447054
rect -1974 443418 -1738 443654
rect -1654 443418 -1418 443654
rect -1974 443098 -1738 443334
rect -1654 443098 -1418 443334
rect 9116 443418 9352 443654
rect 9436 443418 9672 443654
rect 9116 443098 9352 443334
rect 9436 443098 9672 443334
rect 56652 443418 56888 443654
rect 56972 443418 57208 443654
rect 56652 443098 56888 443334
rect 56972 443098 57208 443334
rect 61342 443418 61578 443654
rect 61342 443098 61578 443334
rect 158378 443418 158614 443654
rect 158378 443098 158614 443334
rect 164652 443418 164888 443654
rect 164972 443418 165208 443654
rect 164652 443098 164888 443334
rect 164972 443098 165208 443334
rect 186342 443418 186578 443654
rect 186342 443098 186578 443334
rect 283378 443418 283614 443654
rect 283378 443098 283614 443334
rect 308652 443418 308888 443654
rect 308972 443418 309208 443654
rect 308652 443098 308888 443334
rect 308972 443098 309208 443334
rect 311342 443418 311578 443654
rect 311342 443098 311578 443334
rect 408378 443418 408614 443654
rect 408378 443098 408614 443334
rect 416652 443418 416888 443654
rect 416972 443418 417208 443654
rect 416652 443098 416888 443334
rect 416972 443098 417208 443334
rect 437342 443418 437578 443654
rect 437342 443098 437578 443334
rect 534378 443418 534614 443654
rect 534378 443098 534614 443334
rect 560652 443418 560888 443654
rect 560972 443418 561208 443654
rect 560652 443098 560888 443334
rect 560972 443098 561208 443334
rect 570292 443418 570528 443654
rect 570612 443418 570848 443654
rect 570292 443098 570528 443334
rect 570612 443098 570848 443334
rect 61342 433008 61578 433244
rect 63008 433008 63244 433244
rect 281712 433008 281948 433244
rect 283378 433008 283614 433244
rect 311342 433008 311578 433244
rect 313008 433008 313244 433244
rect 532712 433008 532948 433244
rect 534378 433008 534614 433244
rect 157392 432328 157628 432564
rect 159098 432328 159334 432564
rect 185622 432328 185858 432564
rect 187328 432328 187564 432564
rect 407392 432328 407628 432564
rect 409098 432328 409334 432564
rect 436622 432328 436858 432564
rect 438328 432328 438564 432564
rect 580626 422018 580862 422254
rect 580946 422018 581182 422254
rect 580626 421698 580862 421934
rect 580946 421698 581182 421934
rect 7876 407138 8112 407374
rect 8196 407138 8432 407374
rect 7876 406818 8112 407054
rect 8196 406818 8432 407054
rect 38032 407138 38268 407374
rect 38352 407138 38588 407374
rect 38032 406818 38268 407054
rect 38352 406818 38588 407054
rect 74032 407138 74268 407374
rect 74352 407138 74588 407374
rect 74032 406818 74268 407054
rect 74352 406818 74588 407054
rect 110032 407138 110268 407374
rect 110352 407138 110588 407374
rect 110032 406818 110268 407054
rect 110352 406818 110588 407054
rect 146032 407138 146268 407374
rect 146352 407138 146588 407374
rect 146032 406818 146268 407054
rect 146352 406818 146588 407054
rect 182032 407138 182268 407374
rect 182352 407138 182588 407374
rect 182032 406818 182268 407054
rect 182352 406818 182588 407054
rect 218032 407138 218268 407374
rect 218352 407138 218588 407374
rect 218032 406818 218268 407054
rect 218352 406818 218588 407054
rect 254032 407138 254268 407374
rect 254352 407138 254588 407374
rect 254032 406818 254268 407054
rect 254352 406818 254588 407054
rect 290032 407138 290268 407374
rect 290352 407138 290588 407374
rect 290032 406818 290268 407054
rect 290352 406818 290588 407054
rect 326032 407138 326268 407374
rect 326352 407138 326588 407374
rect 326032 406818 326268 407054
rect 326352 406818 326588 407054
rect 362032 407138 362268 407374
rect 362352 407138 362588 407374
rect 362032 406818 362268 407054
rect 362352 406818 362588 407054
rect 398032 407138 398268 407374
rect 398352 407138 398588 407374
rect 398032 406818 398268 407054
rect 398352 406818 398588 407054
rect 434032 407138 434268 407374
rect 434352 407138 434588 407374
rect 434032 406818 434268 407054
rect 434352 406818 434588 407054
rect 470032 407138 470268 407374
rect 470352 407138 470588 407374
rect 470032 406818 470268 407054
rect 470352 406818 470588 407054
rect 506032 407138 506268 407374
rect 506352 407138 506588 407374
rect 506032 406818 506268 407054
rect 506352 406818 506588 407054
rect 542032 407138 542268 407374
rect 542352 407138 542588 407374
rect 542032 406818 542268 407054
rect 542352 406818 542588 407054
rect 571532 407138 571768 407374
rect 571852 407138 572088 407374
rect 571532 406818 571768 407054
rect 571852 406818 572088 407054
rect -1974 403418 -1738 403654
rect -1654 403418 -1418 403654
rect -1974 403098 -1738 403334
rect -1654 403098 -1418 403334
rect 9116 403418 9352 403654
rect 9436 403418 9672 403654
rect 9116 403098 9352 403334
rect 9436 403098 9672 403334
rect 56652 403418 56888 403654
rect 56972 403418 57208 403654
rect 56652 403098 56888 403334
rect 56972 403098 57208 403334
rect 92652 403418 92888 403654
rect 92972 403418 93208 403654
rect 92652 403098 92888 403334
rect 92972 403098 93208 403334
rect 128652 403418 128888 403654
rect 128972 403418 129208 403654
rect 128652 403098 128888 403334
rect 128972 403098 129208 403334
rect 164652 403418 164888 403654
rect 164972 403418 165208 403654
rect 164652 403098 164888 403334
rect 164972 403098 165208 403334
rect 200652 403418 200888 403654
rect 200972 403418 201208 403654
rect 200652 403098 200888 403334
rect 200972 403098 201208 403334
rect 236652 403418 236888 403654
rect 236972 403418 237208 403654
rect 236652 403098 236888 403334
rect 236972 403098 237208 403334
rect 272652 403418 272888 403654
rect 272972 403418 273208 403654
rect 272652 403098 272888 403334
rect 272972 403098 273208 403334
rect 308652 403418 308888 403654
rect 308972 403418 309208 403654
rect 308652 403098 308888 403334
rect 308972 403098 309208 403334
rect 344652 403418 344888 403654
rect 344972 403418 345208 403654
rect 344652 403098 344888 403334
rect 344972 403098 345208 403334
rect 380652 403418 380888 403654
rect 380972 403418 381208 403654
rect 380652 403098 380888 403334
rect 380972 403098 381208 403334
rect 416652 403418 416888 403654
rect 416972 403418 417208 403654
rect 416652 403098 416888 403334
rect 416972 403098 417208 403334
rect 452652 403418 452888 403654
rect 452972 403418 453208 403654
rect 452652 403098 452888 403334
rect 452972 403098 453208 403334
rect 488652 403418 488888 403654
rect 488972 403418 489208 403654
rect 488652 403098 488888 403334
rect 488972 403098 489208 403334
rect 524652 403418 524888 403654
rect 524972 403418 525208 403654
rect 524652 403098 524888 403334
rect 524972 403098 525208 403334
rect 560652 403418 560888 403654
rect 560972 403418 561208 403654
rect 560652 403098 560888 403334
rect 560972 403098 561208 403334
rect 570292 403418 570528 403654
rect 570612 403418 570848 403654
rect 570292 403098 570528 403334
rect 570612 403098 570848 403334
rect 580626 382018 580862 382254
rect 580946 382018 581182 382254
rect 580626 381698 580862 381934
rect 580946 381698 581182 381934
rect 7876 367138 8112 367374
rect 8196 367138 8432 367374
rect 7876 366818 8112 367054
rect 8196 366818 8432 367054
rect 38032 367138 38268 367374
rect 38352 367138 38588 367374
rect 38032 366818 38268 367054
rect 38352 366818 38588 367054
rect 74032 367138 74268 367374
rect 74352 367138 74588 367374
rect 74032 366818 74268 367054
rect 74352 366818 74588 367054
rect 110032 367138 110268 367374
rect 110352 367138 110588 367374
rect 110032 366818 110268 367054
rect 110352 366818 110588 367054
rect 146032 367138 146268 367374
rect 146352 367138 146588 367374
rect 146032 366818 146268 367054
rect 146352 366818 146588 367054
rect 182032 367138 182268 367374
rect 182352 367138 182588 367374
rect 182032 366818 182268 367054
rect 182352 366818 182588 367054
rect 218032 367138 218268 367374
rect 218352 367138 218588 367374
rect 218032 366818 218268 367054
rect 218352 366818 218588 367054
rect 254032 367138 254268 367374
rect 254352 367138 254588 367374
rect 254032 366818 254268 367054
rect 254352 366818 254588 367054
rect 290032 367138 290268 367374
rect 290352 367138 290588 367374
rect 290032 366818 290268 367054
rect 290352 366818 290588 367054
rect 326032 367138 326268 367374
rect 326352 367138 326588 367374
rect 326032 366818 326268 367054
rect 326352 366818 326588 367054
rect 362032 367138 362268 367374
rect 362352 367138 362588 367374
rect 362032 366818 362268 367054
rect 362352 366818 362588 367054
rect 398032 367138 398268 367374
rect 398352 367138 398588 367374
rect 398032 366818 398268 367054
rect 398352 366818 398588 367054
rect 434032 367138 434268 367374
rect 434352 367138 434588 367374
rect 434032 366818 434268 367054
rect 434352 366818 434588 367054
rect 470032 367138 470268 367374
rect 470352 367138 470588 367374
rect 470032 366818 470268 367054
rect 470352 366818 470588 367054
rect 506032 367138 506268 367374
rect 506352 367138 506588 367374
rect 506032 366818 506268 367054
rect 506352 366818 506588 367054
rect 542032 367138 542268 367374
rect 542352 367138 542588 367374
rect 542032 366818 542268 367054
rect 542352 366818 542588 367054
rect 571532 367138 571768 367374
rect 571852 367138 572088 367374
rect 571532 366818 571768 367054
rect 571852 366818 572088 367054
rect -1974 363418 -1738 363654
rect -1654 363418 -1418 363654
rect -1974 363098 -1738 363334
rect -1654 363098 -1418 363334
rect 9116 363418 9352 363654
rect 9436 363418 9672 363654
rect 9116 363098 9352 363334
rect 9436 363098 9672 363334
rect 56652 363418 56888 363654
rect 56972 363418 57208 363654
rect 56652 363098 56888 363334
rect 56972 363098 57208 363334
rect 92652 363418 92888 363654
rect 92972 363418 93208 363654
rect 92652 363098 92888 363334
rect 92972 363098 93208 363334
rect 128652 363418 128888 363654
rect 128972 363418 129208 363654
rect 128652 363098 128888 363334
rect 128972 363098 129208 363334
rect 164652 363418 164888 363654
rect 164972 363418 165208 363654
rect 164652 363098 164888 363334
rect 164972 363098 165208 363334
rect 200652 363418 200888 363654
rect 200972 363418 201208 363654
rect 200652 363098 200888 363334
rect 200972 363098 201208 363334
rect 236652 363418 236888 363654
rect 236972 363418 237208 363654
rect 236652 363098 236888 363334
rect 236972 363098 237208 363334
rect 272652 363418 272888 363654
rect 272972 363418 273208 363654
rect 272652 363098 272888 363334
rect 272972 363098 273208 363334
rect 308652 363418 308888 363654
rect 308972 363418 309208 363654
rect 308652 363098 308888 363334
rect 308972 363098 309208 363334
rect 344652 363418 344888 363654
rect 344972 363418 345208 363654
rect 344652 363098 344888 363334
rect 344972 363098 345208 363334
rect 380652 363418 380888 363654
rect 380972 363418 381208 363654
rect 380652 363098 380888 363334
rect 380972 363098 381208 363334
rect 416652 363418 416888 363654
rect 416972 363418 417208 363654
rect 416652 363098 416888 363334
rect 416972 363098 417208 363334
rect 452652 363418 452888 363654
rect 452972 363418 453208 363654
rect 452652 363098 452888 363334
rect 452972 363098 453208 363334
rect 488652 363418 488888 363654
rect 488972 363418 489208 363654
rect 488652 363098 488888 363334
rect 488972 363098 489208 363334
rect 524652 363418 524888 363654
rect 524972 363418 525208 363654
rect 524652 363098 524888 363334
rect 524972 363098 525208 363334
rect 560652 363418 560888 363654
rect 560972 363418 561208 363654
rect 560652 363098 560888 363334
rect 560972 363098 561208 363334
rect 570292 363418 570528 363654
rect 570612 363418 570848 363654
rect 570292 363098 570528 363334
rect 570612 363098 570848 363334
rect 580626 342018 580862 342254
rect 580946 342018 581182 342254
rect 580626 341698 580862 341934
rect 580946 341698 581182 341934
rect 7876 327138 8112 327374
rect 8196 327138 8432 327374
rect 7876 326818 8112 327054
rect 8196 326818 8432 327054
rect 38032 327138 38268 327374
rect 38352 327138 38588 327374
rect 38032 326818 38268 327054
rect 38352 326818 38588 327054
rect 74032 327138 74268 327374
rect 74352 327138 74588 327374
rect 74032 326818 74268 327054
rect 74352 326818 74588 327054
rect 110032 327138 110268 327374
rect 110352 327138 110588 327374
rect 110032 326818 110268 327054
rect 110352 326818 110588 327054
rect 146032 327138 146268 327374
rect 146352 327138 146588 327374
rect 146032 326818 146268 327054
rect 146352 326818 146588 327054
rect 182032 327138 182268 327374
rect 182352 327138 182588 327374
rect 182032 326818 182268 327054
rect 182352 326818 182588 327054
rect 218032 327138 218268 327374
rect 218352 327138 218588 327374
rect 218032 326818 218268 327054
rect 218352 326818 218588 327054
rect 254032 327138 254268 327374
rect 254352 327138 254588 327374
rect 254032 326818 254268 327054
rect 254352 326818 254588 327054
rect 290032 327138 290268 327374
rect 290352 327138 290588 327374
rect 290032 326818 290268 327054
rect 290352 326818 290588 327054
rect 326032 327138 326268 327374
rect 326352 327138 326588 327374
rect 326032 326818 326268 327054
rect 326352 326818 326588 327054
rect 362032 327138 362268 327374
rect 362352 327138 362588 327374
rect 362032 326818 362268 327054
rect 362352 326818 362588 327054
rect 398032 327138 398268 327374
rect 398352 327138 398588 327374
rect 398032 326818 398268 327054
rect 398352 326818 398588 327054
rect 434032 327138 434268 327374
rect 434352 327138 434588 327374
rect 434032 326818 434268 327054
rect 434352 326818 434588 327054
rect 470032 327138 470268 327374
rect 470352 327138 470588 327374
rect 470032 326818 470268 327054
rect 470352 326818 470588 327054
rect 506032 327138 506268 327374
rect 506352 327138 506588 327374
rect 506032 326818 506268 327054
rect 506352 326818 506588 327054
rect 542032 327138 542268 327374
rect 542352 327138 542588 327374
rect 542032 326818 542268 327054
rect 542352 326818 542588 327054
rect 571532 327138 571768 327374
rect 571852 327138 572088 327374
rect 571532 326818 571768 327054
rect 571852 326818 572088 327054
rect -1974 323418 -1738 323654
rect -1654 323418 -1418 323654
rect -1974 323098 -1738 323334
rect -1654 323098 -1418 323334
rect 9116 323418 9352 323654
rect 9436 323418 9672 323654
rect 9116 323098 9352 323334
rect 9436 323098 9672 323334
rect 56652 323418 56888 323654
rect 56972 323418 57208 323654
rect 56652 323098 56888 323334
rect 56972 323098 57208 323334
rect 92652 323418 92888 323654
rect 92972 323418 93208 323654
rect 92652 323098 92888 323334
rect 92972 323098 93208 323334
rect 128652 323418 128888 323654
rect 128972 323418 129208 323654
rect 128652 323098 128888 323334
rect 128972 323098 129208 323334
rect 164652 323418 164888 323654
rect 164972 323418 165208 323654
rect 164652 323098 164888 323334
rect 164972 323098 165208 323334
rect 200652 323418 200888 323654
rect 200972 323418 201208 323654
rect 200652 323098 200888 323334
rect 200972 323098 201208 323334
rect 236652 323418 236888 323654
rect 236972 323418 237208 323654
rect 236652 323098 236888 323334
rect 236972 323098 237208 323334
rect 272652 323418 272888 323654
rect 272972 323418 273208 323654
rect 272652 323098 272888 323334
rect 272972 323098 273208 323334
rect 308652 323418 308888 323654
rect 308972 323418 309208 323654
rect 308652 323098 308888 323334
rect 308972 323098 309208 323334
rect 344652 323418 344888 323654
rect 344972 323418 345208 323654
rect 344652 323098 344888 323334
rect 344972 323098 345208 323334
rect 380652 323418 380888 323654
rect 380972 323418 381208 323654
rect 380652 323098 380888 323334
rect 380972 323098 381208 323334
rect 416652 323418 416888 323654
rect 416972 323418 417208 323654
rect 416652 323098 416888 323334
rect 416972 323098 417208 323334
rect 452652 323418 452888 323654
rect 452972 323418 453208 323654
rect 452652 323098 452888 323334
rect 452972 323098 453208 323334
rect 488652 323418 488888 323654
rect 488972 323418 489208 323654
rect 488652 323098 488888 323334
rect 488972 323098 489208 323334
rect 524652 323418 524888 323654
rect 524972 323418 525208 323654
rect 524652 323098 524888 323334
rect 524972 323098 525208 323334
rect 560652 323418 560888 323654
rect 560972 323418 561208 323654
rect 560652 323098 560888 323334
rect 560972 323098 561208 323334
rect 570292 323418 570528 323654
rect 570612 323418 570848 323654
rect 570292 323098 570528 323334
rect 570612 323098 570848 323334
rect 580626 302018 580862 302254
rect 580946 302018 581182 302254
rect 580626 301698 580862 301934
rect 580946 301698 581182 301934
rect 7876 287138 8112 287374
rect 8196 287138 8432 287374
rect 7876 286818 8112 287054
rect 8196 286818 8432 287054
rect 38032 287138 38268 287374
rect 38352 287138 38588 287374
rect 38032 286818 38268 287054
rect 38352 286818 38588 287054
rect 74032 287138 74268 287374
rect 74352 287138 74588 287374
rect 74032 286818 74268 287054
rect 74352 286818 74588 287054
rect 110032 287138 110268 287374
rect 110352 287138 110588 287374
rect 110032 286818 110268 287054
rect 110352 286818 110588 287054
rect 146032 287138 146268 287374
rect 146352 287138 146588 287374
rect 146032 286818 146268 287054
rect 146352 286818 146588 287054
rect 182032 287138 182268 287374
rect 182352 287138 182588 287374
rect 182032 286818 182268 287054
rect 182352 286818 182588 287054
rect 218032 287138 218268 287374
rect 218352 287138 218588 287374
rect 218032 286818 218268 287054
rect 218352 286818 218588 287054
rect 254032 287138 254268 287374
rect 254352 287138 254588 287374
rect 254032 286818 254268 287054
rect 254352 286818 254588 287054
rect 290032 287138 290268 287374
rect 290352 287138 290588 287374
rect 290032 286818 290268 287054
rect 290352 286818 290588 287054
rect 326032 287138 326268 287374
rect 326352 287138 326588 287374
rect 326032 286818 326268 287054
rect 326352 286818 326588 287054
rect 362032 287138 362268 287374
rect 362352 287138 362588 287374
rect 362032 286818 362268 287054
rect 362352 286818 362588 287054
rect 398032 287138 398268 287374
rect 398352 287138 398588 287374
rect 398032 286818 398268 287054
rect 398352 286818 398588 287054
rect 434032 287138 434268 287374
rect 434352 287138 434588 287374
rect 434032 286818 434268 287054
rect 434352 286818 434588 287054
rect 470032 287138 470268 287374
rect 470352 287138 470588 287374
rect 470032 286818 470268 287054
rect 470352 286818 470588 287054
rect 506032 287138 506268 287374
rect 506352 287138 506588 287374
rect 506032 286818 506268 287054
rect 506352 286818 506588 287054
rect 542032 287138 542268 287374
rect 542352 287138 542588 287374
rect 542032 286818 542268 287054
rect 542352 286818 542588 287054
rect 571532 287138 571768 287374
rect 571852 287138 572088 287374
rect 571532 286818 571768 287054
rect 571852 286818 572088 287054
rect -1974 283418 -1738 283654
rect -1654 283418 -1418 283654
rect -1974 283098 -1738 283334
rect -1654 283098 -1418 283334
rect 9116 283418 9352 283654
rect 9436 283418 9672 283654
rect 9116 283098 9352 283334
rect 9436 283098 9672 283334
rect 56652 283418 56888 283654
rect 56972 283418 57208 283654
rect 56652 283098 56888 283334
rect 56972 283098 57208 283334
rect 92652 283418 92888 283654
rect 92972 283418 93208 283654
rect 92652 283098 92888 283334
rect 92972 283098 93208 283334
rect 128652 283418 128888 283654
rect 128972 283418 129208 283654
rect 128652 283098 128888 283334
rect 128972 283098 129208 283334
rect 164652 283418 164888 283654
rect 164972 283418 165208 283654
rect 164652 283098 164888 283334
rect 164972 283098 165208 283334
rect 200652 283418 200888 283654
rect 200972 283418 201208 283654
rect 200652 283098 200888 283334
rect 200972 283098 201208 283334
rect 236652 283418 236888 283654
rect 236972 283418 237208 283654
rect 236652 283098 236888 283334
rect 236972 283098 237208 283334
rect 272652 283418 272888 283654
rect 272972 283418 273208 283654
rect 272652 283098 272888 283334
rect 272972 283098 273208 283334
rect 308652 283418 308888 283654
rect 308972 283418 309208 283654
rect 308652 283098 308888 283334
rect 308972 283098 309208 283334
rect 344652 283418 344888 283654
rect 344972 283418 345208 283654
rect 344652 283098 344888 283334
rect 344972 283098 345208 283334
rect 380652 283418 380888 283654
rect 380972 283418 381208 283654
rect 380652 283098 380888 283334
rect 380972 283098 381208 283334
rect 416652 283418 416888 283654
rect 416972 283418 417208 283654
rect 416652 283098 416888 283334
rect 416972 283098 417208 283334
rect 452652 283418 452888 283654
rect 452972 283418 453208 283654
rect 452652 283098 452888 283334
rect 452972 283098 453208 283334
rect 488652 283418 488888 283654
rect 488972 283418 489208 283654
rect 488652 283098 488888 283334
rect 488972 283098 489208 283334
rect 524652 283418 524888 283654
rect 524972 283418 525208 283654
rect 524652 283098 524888 283334
rect 524972 283098 525208 283334
rect 560652 283418 560888 283654
rect 560972 283418 561208 283654
rect 560652 283098 560888 283334
rect 560972 283098 561208 283334
rect 570292 283418 570528 283654
rect 570612 283418 570848 283654
rect 570292 283098 570528 283334
rect 570612 283098 570848 283334
rect 580626 262018 580862 262254
rect 580946 262018 581182 262254
rect 580626 261698 580862 261934
rect 580946 261698 581182 261934
rect 7876 247138 8112 247374
rect 8196 247138 8432 247374
rect 7876 246818 8112 247054
rect 8196 246818 8432 247054
rect 38032 247138 38268 247374
rect 38352 247138 38588 247374
rect 38032 246818 38268 247054
rect 38352 246818 38588 247054
rect 74032 247138 74268 247374
rect 74352 247138 74588 247374
rect 74032 246818 74268 247054
rect 74352 246818 74588 247054
rect 110032 247138 110268 247374
rect 110352 247138 110588 247374
rect 110032 246818 110268 247054
rect 110352 246818 110588 247054
rect 146032 247138 146268 247374
rect 146352 247138 146588 247374
rect 146032 246818 146268 247054
rect 146352 246818 146588 247054
rect 182032 247138 182268 247374
rect 182352 247138 182588 247374
rect 182032 246818 182268 247054
rect 182352 246818 182588 247054
rect 218032 247138 218268 247374
rect 218352 247138 218588 247374
rect 218032 246818 218268 247054
rect 218352 246818 218588 247054
rect 254032 247138 254268 247374
rect 254352 247138 254588 247374
rect 254032 246818 254268 247054
rect 254352 246818 254588 247054
rect 290032 247138 290268 247374
rect 290352 247138 290588 247374
rect 290032 246818 290268 247054
rect 290352 246818 290588 247054
rect 326032 247138 326268 247374
rect 326352 247138 326588 247374
rect 326032 246818 326268 247054
rect 326352 246818 326588 247054
rect 362032 247138 362268 247374
rect 362352 247138 362588 247374
rect 362032 246818 362268 247054
rect 362352 246818 362588 247054
rect 398032 247138 398268 247374
rect 398352 247138 398588 247374
rect 398032 246818 398268 247054
rect 398352 246818 398588 247054
rect 434032 247138 434268 247374
rect 434352 247138 434588 247374
rect 434032 246818 434268 247054
rect 434352 246818 434588 247054
rect 470032 247138 470268 247374
rect 470352 247138 470588 247374
rect 470032 246818 470268 247054
rect 470352 246818 470588 247054
rect 506032 247138 506268 247374
rect 506352 247138 506588 247374
rect 506032 246818 506268 247054
rect 506352 246818 506588 247054
rect 542032 247138 542268 247374
rect 542352 247138 542588 247374
rect 542032 246818 542268 247054
rect 542352 246818 542588 247054
rect 571532 247138 571768 247374
rect 571852 247138 572088 247374
rect 571532 246818 571768 247054
rect 571852 246818 572088 247054
rect -1974 243418 -1738 243654
rect -1654 243418 -1418 243654
rect -1974 243098 -1738 243334
rect -1654 243098 -1418 243334
rect 9116 243418 9352 243654
rect 9436 243418 9672 243654
rect 9116 243098 9352 243334
rect 9436 243098 9672 243334
rect 56652 243418 56888 243654
rect 56972 243418 57208 243654
rect 56652 243098 56888 243334
rect 56972 243098 57208 243334
rect 92652 243418 92888 243654
rect 92972 243418 93208 243654
rect 92652 243098 92888 243334
rect 92972 243098 93208 243334
rect 128652 243418 128888 243654
rect 128972 243418 129208 243654
rect 128652 243098 128888 243334
rect 128972 243098 129208 243334
rect 164652 243418 164888 243654
rect 164972 243418 165208 243654
rect 164652 243098 164888 243334
rect 164972 243098 165208 243334
rect 200652 243418 200888 243654
rect 200972 243418 201208 243654
rect 200652 243098 200888 243334
rect 200972 243098 201208 243334
rect 236652 243418 236888 243654
rect 236972 243418 237208 243654
rect 236652 243098 236888 243334
rect 236972 243098 237208 243334
rect 272652 243418 272888 243654
rect 272972 243418 273208 243654
rect 272652 243098 272888 243334
rect 272972 243098 273208 243334
rect 308652 243418 308888 243654
rect 308972 243418 309208 243654
rect 308652 243098 308888 243334
rect 308972 243098 309208 243334
rect 344652 243418 344888 243654
rect 344972 243418 345208 243654
rect 344652 243098 344888 243334
rect 344972 243098 345208 243334
rect 380652 243418 380888 243654
rect 380972 243418 381208 243654
rect 380652 243098 380888 243334
rect 380972 243098 381208 243334
rect 416652 243418 416888 243654
rect 416972 243418 417208 243654
rect 416652 243098 416888 243334
rect 416972 243098 417208 243334
rect 452652 243418 452888 243654
rect 452972 243418 453208 243654
rect 452652 243098 452888 243334
rect 452972 243098 453208 243334
rect 488652 243418 488888 243654
rect 488972 243418 489208 243654
rect 488652 243098 488888 243334
rect 488972 243098 489208 243334
rect 524652 243418 524888 243654
rect 524972 243418 525208 243654
rect 524652 243098 524888 243334
rect 524972 243098 525208 243334
rect 560652 243418 560888 243654
rect 560972 243418 561208 243654
rect 560652 243098 560888 243334
rect 560972 243098 561208 243334
rect 570292 243418 570528 243654
rect 570612 243418 570848 243654
rect 570292 243098 570528 243334
rect 570612 243098 570848 243334
rect 580626 222018 580862 222254
rect 580946 222018 581182 222254
rect 580626 221698 580862 221934
rect 580946 221698 581182 221934
rect 7876 207138 8112 207374
rect 8196 207138 8432 207374
rect 7876 206818 8112 207054
rect 8196 206818 8432 207054
rect 38032 207138 38268 207374
rect 38352 207138 38588 207374
rect 38032 206818 38268 207054
rect 38352 206818 38588 207054
rect 74032 207138 74268 207374
rect 74352 207138 74588 207374
rect 74032 206818 74268 207054
rect 74352 206818 74588 207054
rect 110032 207138 110268 207374
rect 110352 207138 110588 207374
rect 110032 206818 110268 207054
rect 110352 206818 110588 207054
rect 146032 207138 146268 207374
rect 146352 207138 146588 207374
rect 146032 206818 146268 207054
rect 146352 206818 146588 207054
rect 182032 207138 182268 207374
rect 182352 207138 182588 207374
rect 182032 206818 182268 207054
rect 182352 206818 182588 207054
rect 218032 207138 218268 207374
rect 218352 207138 218588 207374
rect 218032 206818 218268 207054
rect 218352 206818 218588 207054
rect 254032 207138 254268 207374
rect 254352 207138 254588 207374
rect 254032 206818 254268 207054
rect 254352 206818 254588 207054
rect 290032 207138 290268 207374
rect 290352 207138 290588 207374
rect 290032 206818 290268 207054
rect 290352 206818 290588 207054
rect 326032 207138 326268 207374
rect 326352 207138 326588 207374
rect 326032 206818 326268 207054
rect 326352 206818 326588 207054
rect 362032 207138 362268 207374
rect 362352 207138 362588 207374
rect 362032 206818 362268 207054
rect 362352 206818 362588 207054
rect 398032 207138 398268 207374
rect 398352 207138 398588 207374
rect 398032 206818 398268 207054
rect 398352 206818 398588 207054
rect 434032 207138 434268 207374
rect 434352 207138 434588 207374
rect 434032 206818 434268 207054
rect 434352 206818 434588 207054
rect 470032 207138 470268 207374
rect 470352 207138 470588 207374
rect 470032 206818 470268 207054
rect 470352 206818 470588 207054
rect 506032 207138 506268 207374
rect 506352 207138 506588 207374
rect 506032 206818 506268 207054
rect 506352 206818 506588 207054
rect 542032 207138 542268 207374
rect 542352 207138 542588 207374
rect 542032 206818 542268 207054
rect 542352 206818 542588 207054
rect 571532 207138 571768 207374
rect 571852 207138 572088 207374
rect 571532 206818 571768 207054
rect 571852 206818 572088 207054
rect -1974 203418 -1738 203654
rect -1654 203418 -1418 203654
rect -1974 203098 -1738 203334
rect -1654 203098 -1418 203334
rect 9116 203418 9352 203654
rect 9436 203418 9672 203654
rect 9116 203098 9352 203334
rect 9436 203098 9672 203334
rect 56652 203418 56888 203654
rect 56972 203418 57208 203654
rect 56652 203098 56888 203334
rect 56972 203098 57208 203334
rect 92652 203418 92888 203654
rect 92972 203418 93208 203654
rect 92652 203098 92888 203334
rect 92972 203098 93208 203334
rect 128652 203418 128888 203654
rect 128972 203418 129208 203654
rect 128652 203098 128888 203334
rect 128972 203098 129208 203334
rect 164652 203418 164888 203654
rect 164972 203418 165208 203654
rect 164652 203098 164888 203334
rect 164972 203098 165208 203334
rect 200652 203418 200888 203654
rect 200972 203418 201208 203654
rect 200652 203098 200888 203334
rect 200972 203098 201208 203334
rect 236652 203418 236888 203654
rect 236972 203418 237208 203654
rect 236652 203098 236888 203334
rect 236972 203098 237208 203334
rect 272652 203418 272888 203654
rect 272972 203418 273208 203654
rect 272652 203098 272888 203334
rect 272972 203098 273208 203334
rect 308652 203418 308888 203654
rect 308972 203418 309208 203654
rect 308652 203098 308888 203334
rect 308972 203098 309208 203334
rect 344652 203418 344888 203654
rect 344972 203418 345208 203654
rect 344652 203098 344888 203334
rect 344972 203098 345208 203334
rect 380652 203418 380888 203654
rect 380972 203418 381208 203654
rect 380652 203098 380888 203334
rect 380972 203098 381208 203334
rect 416652 203418 416888 203654
rect 416972 203418 417208 203654
rect 416652 203098 416888 203334
rect 416972 203098 417208 203334
rect 452652 203418 452888 203654
rect 452972 203418 453208 203654
rect 452652 203098 452888 203334
rect 452972 203098 453208 203334
rect 488652 203418 488888 203654
rect 488972 203418 489208 203654
rect 488652 203098 488888 203334
rect 488972 203098 489208 203334
rect 524652 203418 524888 203654
rect 524972 203418 525208 203654
rect 524652 203098 524888 203334
rect 524972 203098 525208 203334
rect 560652 203418 560888 203654
rect 560972 203418 561208 203654
rect 560652 203098 560888 203334
rect 560972 203098 561208 203334
rect 570292 203418 570528 203654
rect 570612 203418 570848 203654
rect 570292 203098 570528 203334
rect 570612 203098 570848 203334
rect 580626 182018 580862 182254
rect 580946 182018 581182 182254
rect 580626 181698 580862 181934
rect 580946 181698 581182 181934
rect 7876 167138 8112 167374
rect 8196 167138 8432 167374
rect 7876 166818 8112 167054
rect 8196 166818 8432 167054
rect 38032 167138 38268 167374
rect 38352 167138 38588 167374
rect 38032 166818 38268 167054
rect 38352 166818 38588 167054
rect 60622 167138 60858 167374
rect 60622 166818 60858 167054
rect 159098 167138 159334 167374
rect 159098 166818 159334 167054
rect 182032 167138 182268 167374
rect 182352 167138 182588 167374
rect 182032 166818 182268 167054
rect 182352 166818 182588 167054
rect 185622 167138 185858 167374
rect 185622 166818 185858 167054
rect 284098 167138 284334 167374
rect 284098 166818 284334 167054
rect 290032 167138 290268 167374
rect 290352 167138 290588 167374
rect 290032 166818 290268 167054
rect 290352 166818 290588 167054
rect 310622 167138 310858 167374
rect 310622 166818 310858 167054
rect 409098 167138 409334 167374
rect 409098 166818 409334 167054
rect 434032 167138 434268 167374
rect 434352 167138 434588 167374
rect 434032 166818 434268 167054
rect 434352 166818 434588 167054
rect 436622 167138 436858 167374
rect 436622 166818 436858 167054
rect 535098 167138 535334 167374
rect 535098 166818 535334 167054
rect 542032 167138 542268 167374
rect 542352 167138 542588 167374
rect 542032 166818 542268 167054
rect 542352 166818 542588 167054
rect 571532 167138 571768 167374
rect 571852 167138 572088 167374
rect 571532 166818 571768 167054
rect 571852 166818 572088 167054
rect -1974 163418 -1738 163654
rect -1654 163418 -1418 163654
rect -1974 163098 -1738 163334
rect -1654 163098 -1418 163334
rect 9116 163418 9352 163654
rect 9436 163418 9672 163654
rect 9116 163098 9352 163334
rect 9436 163098 9672 163334
rect 56652 163418 56888 163654
rect 56972 163418 57208 163654
rect 56652 163098 56888 163334
rect 56972 163098 57208 163334
rect 61342 163418 61578 163654
rect 61342 163098 61578 163334
rect 158378 163418 158614 163654
rect 158378 163098 158614 163334
rect 164652 163418 164888 163654
rect 164972 163418 165208 163654
rect 164652 163098 164888 163334
rect 164972 163098 165208 163334
rect 186342 163418 186578 163654
rect 186342 163098 186578 163334
rect 283378 163418 283614 163654
rect 283378 163098 283614 163334
rect 308652 163418 308888 163654
rect 308972 163418 309208 163654
rect 308652 163098 308888 163334
rect 308972 163098 309208 163334
rect 311342 163418 311578 163654
rect 311342 163098 311578 163334
rect 408378 163418 408614 163654
rect 408378 163098 408614 163334
rect 416652 163418 416888 163654
rect 416972 163418 417208 163654
rect 416652 163098 416888 163334
rect 416972 163098 417208 163334
rect 437342 163418 437578 163654
rect 437342 163098 437578 163334
rect 534378 163418 534614 163654
rect 534378 163098 534614 163334
rect 560652 163418 560888 163654
rect 560972 163418 561208 163654
rect 560652 163098 560888 163334
rect 560972 163098 561208 163334
rect 570292 163418 570528 163654
rect 570612 163418 570848 163654
rect 570292 163098 570528 163334
rect 570612 163098 570848 163334
rect 580626 142018 580862 142254
rect 580946 142018 581182 142254
rect 580626 141698 580862 141934
rect 580946 141698 581182 141934
rect 7876 127138 8112 127374
rect 8196 127138 8432 127374
rect 7876 126818 8112 127054
rect 8196 126818 8432 127054
rect 38032 127138 38268 127374
rect 38352 127138 38588 127374
rect 38032 126818 38268 127054
rect 38352 126818 38588 127054
rect 60622 127138 60858 127374
rect 60622 126818 60858 127054
rect 159098 127138 159334 127374
rect 159098 126818 159334 127054
rect 182032 127138 182268 127374
rect 182352 127138 182588 127374
rect 182032 126818 182268 127054
rect 182352 126818 182588 127054
rect 185622 127138 185858 127374
rect 185622 126818 185858 127054
rect 284098 127138 284334 127374
rect 284098 126818 284334 127054
rect 290032 127138 290268 127374
rect 290352 127138 290588 127374
rect 290032 126818 290268 127054
rect 290352 126818 290588 127054
rect 310622 127138 310858 127374
rect 310622 126818 310858 127054
rect 409098 127138 409334 127374
rect 409098 126818 409334 127054
rect 434032 127138 434268 127374
rect 434352 127138 434588 127374
rect 434032 126818 434268 127054
rect 434352 126818 434588 127054
rect 436622 127138 436858 127374
rect 436622 126818 436858 127054
rect 535098 127138 535334 127374
rect 535098 126818 535334 127054
rect 542032 127138 542268 127374
rect 542352 127138 542588 127374
rect 542032 126818 542268 127054
rect 542352 126818 542588 127054
rect 571532 127138 571768 127374
rect 571852 127138 572088 127374
rect 571532 126818 571768 127054
rect 571852 126818 572088 127054
rect -1974 123418 -1738 123654
rect -1654 123418 -1418 123654
rect -1974 123098 -1738 123334
rect -1654 123098 -1418 123334
rect 9116 123418 9352 123654
rect 9436 123418 9672 123654
rect 9116 123098 9352 123334
rect 9436 123098 9672 123334
rect 56652 123418 56888 123654
rect 56972 123418 57208 123654
rect 56652 123098 56888 123334
rect 56972 123098 57208 123334
rect 61342 123418 61578 123654
rect 61342 123098 61578 123334
rect 158378 123418 158614 123654
rect 158378 123098 158614 123334
rect 164652 123418 164888 123654
rect 164972 123418 165208 123654
rect 164652 123098 164888 123334
rect 164972 123098 165208 123334
rect 186342 123418 186578 123654
rect 186342 123098 186578 123334
rect 283378 123418 283614 123654
rect 283378 123098 283614 123334
rect 308652 123418 308888 123654
rect 308972 123418 309208 123654
rect 308652 123098 308888 123334
rect 308972 123098 309208 123334
rect 311342 123418 311578 123654
rect 311342 123098 311578 123334
rect 408378 123418 408614 123654
rect 408378 123098 408614 123334
rect 416652 123418 416888 123654
rect 416972 123418 417208 123654
rect 416652 123098 416888 123334
rect 416972 123098 417208 123334
rect 437342 123418 437578 123654
rect 437342 123098 437578 123334
rect 534378 123418 534614 123654
rect 534378 123098 534614 123334
rect 560652 123418 560888 123654
rect 560972 123418 561208 123654
rect 560652 123098 560888 123334
rect 560972 123098 561208 123334
rect 570292 123418 570528 123654
rect 570612 123418 570848 123654
rect 570292 123098 570528 123334
rect 570612 123098 570848 123334
rect 61342 121008 61578 121244
rect 63008 121008 63244 121244
rect 281712 121008 281948 121244
rect 283378 121008 283614 121244
rect 311342 121008 311578 121244
rect 313008 121008 313244 121244
rect 532712 121008 532948 121244
rect 534378 121008 534614 121244
rect 157392 120328 157628 120564
rect 159098 120328 159334 120564
rect 185622 120328 185858 120564
rect 187328 120328 187564 120564
rect 407392 120328 407628 120564
rect 409098 120328 409334 120564
rect 436622 120328 436858 120564
rect 438328 120328 438564 120564
rect 580626 102018 580862 102254
rect 580946 102018 581182 102254
rect 580626 101698 580862 101934
rect 580946 101698 581182 101934
rect 7876 87138 8112 87374
rect 8196 87138 8432 87374
rect 7876 86818 8112 87054
rect 8196 86818 8432 87054
rect 38032 87138 38268 87374
rect 38352 87138 38588 87374
rect 38032 86818 38268 87054
rect 38352 86818 38588 87054
rect 60622 87138 60858 87374
rect 60622 86818 60858 87054
rect 159098 87138 159334 87374
rect 159098 86818 159334 87054
rect 182032 87138 182268 87374
rect 182352 87138 182588 87374
rect 182032 86818 182268 87054
rect 182352 86818 182588 87054
rect 185622 87138 185858 87374
rect 185622 86818 185858 87054
rect 284098 87138 284334 87374
rect 284098 86818 284334 87054
rect 290032 87138 290268 87374
rect 290352 87138 290588 87374
rect 290032 86818 290268 87054
rect 290352 86818 290588 87054
rect 310622 87138 310858 87374
rect 310622 86818 310858 87054
rect 409098 87138 409334 87374
rect 409098 86818 409334 87054
rect 434032 87138 434268 87374
rect 434352 87138 434588 87374
rect 434032 86818 434268 87054
rect 434352 86818 434588 87054
rect 436622 87138 436858 87374
rect 436622 86818 436858 87054
rect 535098 87138 535334 87374
rect 535098 86818 535334 87054
rect 542032 87138 542268 87374
rect 542352 87138 542588 87374
rect 542032 86818 542268 87054
rect 542352 86818 542588 87054
rect 571532 87138 571768 87374
rect 571852 87138 572088 87374
rect 571532 86818 571768 87054
rect 571852 86818 572088 87054
rect -1974 83418 -1738 83654
rect -1654 83418 -1418 83654
rect -1974 83098 -1738 83334
rect -1654 83098 -1418 83334
rect 9116 83418 9352 83654
rect 9436 83418 9672 83654
rect 9116 83098 9352 83334
rect 9436 83098 9672 83334
rect 56652 83418 56888 83654
rect 56972 83418 57208 83654
rect 56652 83098 56888 83334
rect 56972 83098 57208 83334
rect 61342 83418 61578 83654
rect 61342 83098 61578 83334
rect 158378 83418 158614 83654
rect 158378 83098 158614 83334
rect 164652 83418 164888 83654
rect 164972 83418 165208 83654
rect 164652 83098 164888 83334
rect 164972 83098 165208 83334
rect 186342 83418 186578 83654
rect 186342 83098 186578 83334
rect 283378 83418 283614 83654
rect 283378 83098 283614 83334
rect 308652 83418 308888 83654
rect 308972 83418 309208 83654
rect 308652 83098 308888 83334
rect 308972 83098 309208 83334
rect 311342 83418 311578 83654
rect 311342 83098 311578 83334
rect 408378 83418 408614 83654
rect 408378 83098 408614 83334
rect 416652 83418 416888 83654
rect 416972 83418 417208 83654
rect 416652 83098 416888 83334
rect 416972 83098 417208 83334
rect 437342 83418 437578 83654
rect 437342 83098 437578 83334
rect 534378 83418 534614 83654
rect 534378 83098 534614 83334
rect 560652 83418 560888 83654
rect 560972 83418 561208 83654
rect 560652 83098 560888 83334
rect 560972 83098 561208 83334
rect 570292 83418 570528 83654
rect 570612 83418 570848 83654
rect 570292 83098 570528 83334
rect 570612 83098 570848 83334
rect 580626 62018 580862 62254
rect 580946 62018 581182 62254
rect 580626 61698 580862 61934
rect 580946 61698 581182 61934
rect 7876 47138 8112 47374
rect 8196 47138 8432 47374
rect 7876 46818 8112 47054
rect 8196 46818 8432 47054
rect 38032 47138 38268 47374
rect 38352 47138 38588 47374
rect 38032 46818 38268 47054
rect 38352 46818 38588 47054
rect 60622 47138 60858 47374
rect 60622 46818 60858 47054
rect 159098 47138 159334 47374
rect 159098 46818 159334 47054
rect 182032 47138 182268 47374
rect 182352 47138 182588 47374
rect 182032 46818 182268 47054
rect 182352 46818 182588 47054
rect 185622 47138 185858 47374
rect 185622 46818 185858 47054
rect 284098 47138 284334 47374
rect 284098 46818 284334 47054
rect 290032 47138 290268 47374
rect 290352 47138 290588 47374
rect 290032 46818 290268 47054
rect 290352 46818 290588 47054
rect 310622 47138 310858 47374
rect 310622 46818 310858 47054
rect 409098 47138 409334 47374
rect 409098 46818 409334 47054
rect 434032 47138 434268 47374
rect 434352 47138 434588 47374
rect 434032 46818 434268 47054
rect 434352 46818 434588 47054
rect 436622 47138 436858 47374
rect 436622 46818 436858 47054
rect 535098 47138 535334 47374
rect 535098 46818 535334 47054
rect 542032 47138 542268 47374
rect 542352 47138 542588 47374
rect 542032 46818 542268 47054
rect 542352 46818 542588 47054
rect 571532 47138 571768 47374
rect 571852 47138 572088 47374
rect 571532 46818 571768 47054
rect 571852 46818 572088 47054
rect -1974 43418 -1738 43654
rect -1654 43418 -1418 43654
rect -1974 43098 -1738 43334
rect -1654 43098 -1418 43334
rect 9116 43418 9352 43654
rect 9436 43418 9672 43654
rect 9116 43098 9352 43334
rect 9436 43098 9672 43334
rect 56652 43418 56888 43654
rect 56972 43418 57208 43654
rect 56652 43098 56888 43334
rect 56972 43098 57208 43334
rect 61342 43418 61578 43654
rect 61342 43098 61578 43334
rect 158378 43418 158614 43654
rect 158378 43098 158614 43334
rect 164652 43418 164888 43654
rect 164972 43418 165208 43654
rect 164652 43098 164888 43334
rect 164972 43098 165208 43334
rect 186342 43418 186578 43654
rect 186342 43098 186578 43334
rect 283378 43418 283614 43654
rect 283378 43098 283614 43334
rect 308652 43418 308888 43654
rect 308972 43418 309208 43654
rect 308652 43098 308888 43334
rect 308972 43098 309208 43334
rect 311342 43418 311578 43654
rect 311342 43098 311578 43334
rect 408378 43418 408614 43654
rect 408378 43098 408614 43334
rect 416652 43418 416888 43654
rect 416972 43418 417208 43654
rect 416652 43098 416888 43334
rect 416972 43098 417208 43334
rect 437342 43418 437578 43654
rect 437342 43098 437578 43334
rect 534378 43418 534614 43654
rect 534378 43098 534614 43334
rect 560652 43418 560888 43654
rect 560972 43418 561208 43654
rect 560652 43098 560888 43334
rect 560972 43098 561208 43334
rect 570292 43418 570528 43654
rect 570612 43418 570848 43654
rect 570292 43098 570528 43334
rect 570612 43098 570848 43334
rect 580626 22018 580862 22254
rect 580946 22018 581182 22254
rect 580626 21698 580862 21934
rect 580946 21698 581182 21934
rect 61342 21008 61578 21244
rect 63008 21008 63244 21244
rect 188008 21008 188244 21244
rect 311342 21008 311578 21244
rect 313008 21008 313244 21244
rect 439008 21008 439244 21244
rect 62328 20328 62564 20564
rect 185622 20328 185858 20564
rect 187328 20328 187564 20564
rect 312328 20328 312564 20564
rect 436622 20328 436858 20564
rect 438328 20328 438564 20564
rect 62328 19598 62564 19834
rect 188008 19342 188244 19578
rect 312328 19598 312564 19834
rect 439008 19342 439244 19578
rect 9116 9444 9352 9680
rect 9436 9444 9672 9680
rect 9116 9124 9352 9360
rect 9436 9124 9672 9360
rect 56652 9444 56888 9680
rect 56972 9444 57208 9680
rect 56652 9124 56888 9360
rect 56972 9124 57208 9360
rect 92652 9444 92888 9680
rect 92972 9444 93208 9680
rect 92652 9124 92888 9360
rect 92972 9124 93208 9360
rect 128652 9444 128888 9680
rect 128972 9444 129208 9680
rect 128652 9124 128888 9360
rect 128972 9124 129208 9360
rect 164652 9444 164888 9680
rect 164972 9444 165208 9680
rect 164652 9124 164888 9360
rect 164972 9124 165208 9360
rect 200652 9444 200888 9680
rect 200972 9444 201208 9680
rect 200652 9124 200888 9360
rect 200972 9124 201208 9360
rect 236652 9444 236888 9680
rect 236972 9444 237208 9680
rect 236652 9124 236888 9360
rect 236972 9124 237208 9360
rect 272652 9444 272888 9680
rect 272972 9444 273208 9680
rect 272652 9124 272888 9360
rect 272972 9124 273208 9360
rect 308652 9444 308888 9680
rect 308972 9444 309208 9680
rect 308652 9124 308888 9360
rect 308972 9124 309208 9360
rect 344652 9444 344888 9680
rect 344972 9444 345208 9680
rect 344652 9124 344888 9360
rect 344972 9124 345208 9360
rect 380652 9444 380888 9680
rect 380972 9444 381208 9680
rect 380652 9124 380888 9360
rect 380972 9124 381208 9360
rect 416652 9444 416888 9680
rect 416972 9444 417208 9680
rect 416652 9124 416888 9360
rect 416972 9124 417208 9360
rect 452652 9444 452888 9680
rect 452972 9444 453208 9680
rect 452652 9124 452888 9360
rect 452972 9124 453208 9360
rect 488652 9444 488888 9680
rect 488972 9444 489208 9680
rect 488652 9124 488888 9360
rect 488972 9124 489208 9360
rect 524652 9444 524888 9680
rect 524972 9444 525208 9680
rect 524652 9124 524888 9360
rect 524972 9124 525208 9360
rect 560652 9444 560888 9680
rect 560972 9444 561208 9680
rect 560652 9124 560888 9360
rect 560972 9124 561208 9360
rect 570292 9444 570528 9680
rect 570612 9444 570848 9680
rect 570292 9124 570528 9360
rect 570612 9124 570848 9360
rect 7876 8204 8112 8440
rect 8196 8204 8432 8440
rect 7876 7884 8112 8120
rect 8196 7884 8432 8120
rect 38032 8204 38268 8440
rect 38352 8204 38588 8440
rect 38032 7884 38268 8120
rect 38352 7884 38588 8120
rect 74032 8204 74268 8440
rect 74352 8204 74588 8440
rect 74032 7884 74268 8120
rect 74352 7884 74588 8120
rect 110032 8204 110268 8440
rect 110352 8204 110588 8440
rect 110032 7884 110268 8120
rect 110352 7884 110588 8120
rect 146032 8204 146268 8440
rect 146352 8204 146588 8440
rect 146032 7884 146268 8120
rect 146352 7884 146588 8120
rect 182032 8204 182268 8440
rect 182352 8204 182588 8440
rect 182032 7884 182268 8120
rect 182352 7884 182588 8120
rect 218032 8204 218268 8440
rect 218352 8204 218588 8440
rect 218032 7884 218268 8120
rect 218352 7884 218588 8120
rect 254032 8204 254268 8440
rect 254352 8204 254588 8440
rect 254032 7884 254268 8120
rect 254352 7884 254588 8120
rect 290032 8204 290268 8440
rect 290352 8204 290588 8440
rect 290032 7884 290268 8120
rect 290352 7884 290588 8120
rect 326032 8204 326268 8440
rect 326352 8204 326588 8440
rect 326032 7884 326268 8120
rect 326352 7884 326588 8120
rect 362032 8204 362268 8440
rect 362352 8204 362588 8440
rect 362032 7884 362268 8120
rect 362352 7884 362588 8120
rect 398032 8204 398268 8440
rect 398352 8204 398588 8440
rect 398032 7884 398268 8120
rect 398352 7884 398588 8120
rect 434032 8204 434268 8440
rect 434352 8204 434588 8440
rect 434032 7884 434268 8120
rect 434352 7884 434588 8120
rect 470032 8204 470268 8440
rect 470352 8204 470588 8440
rect 470032 7884 470268 8120
rect 470352 7884 470588 8120
rect 506032 8204 506268 8440
rect 506352 8204 506588 8440
rect 506032 7884 506268 8120
rect 506352 7884 506588 8120
rect 542032 8204 542268 8440
rect 542352 8204 542588 8440
rect 542032 7884 542268 8120
rect 542352 7884 542588 8120
rect 571532 8204 571768 8440
rect 571852 8204 572088 8440
rect 571532 7884 571768 8120
rect 571852 7884 572088 8120
rect 7876 7138 8112 7374
rect 8196 7138 8432 7374
rect 7876 6818 8112 7054
rect 8196 6818 8432 7054
rect 571532 7138 571768 7374
rect 571852 7138 572088 7374
rect 571532 6818 571768 7054
rect 571852 6818 572088 7054
rect -1974 3418 -1738 3654
rect -1654 3418 -1418 3654
rect -1974 3098 -1738 3334
rect -1654 3098 -1418 3334
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect -5084 -3692 -4848 -3456
rect -4764 -3692 -4528 -3456
rect -5084 -4012 -4848 -3776
rect -4764 -4012 -4528 -3776
rect -8194 -6802 -7958 -6566
rect -7874 -6802 -7638 -6566
rect -8194 -7122 -7958 -6886
rect -7874 -7122 -7638 -6886
rect -11304 -9912 -11068 -9676
rect -10984 -9912 -10748 -9676
rect -11304 -10232 -11068 -9996
rect -10984 -10232 -10748 -9996
rect -14414 -13022 -14178 -12786
rect -14094 -13022 -13858 -12786
rect -14414 -13342 -14178 -13106
rect -14094 -13342 -13858 -13106
rect -17524 -16132 -17288 -15896
rect -17204 -16132 -16968 -15896
rect -17524 -16452 -17288 -16216
rect -17204 -16452 -16968 -16216
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 683418 585578 683654
rect 585662 683418 585898 683654
rect 585342 683098 585578 683334
rect 585662 683098 585898 683334
rect 585342 643418 585578 643654
rect 585662 643418 585898 643654
rect 585342 643098 585578 643334
rect 585662 643098 585898 643334
rect 585342 603418 585578 603654
rect 585662 603418 585898 603654
rect 585342 603098 585578 603334
rect 585662 603098 585898 603334
rect 585342 563418 585578 563654
rect 585662 563418 585898 563654
rect 585342 563098 585578 563334
rect 585662 563098 585898 563334
rect 585342 523418 585578 523654
rect 585662 523418 585898 523654
rect 585342 523098 585578 523334
rect 585662 523098 585898 523334
rect 585342 483418 585578 483654
rect 585662 483418 585898 483654
rect 585342 483098 585578 483334
rect 585662 483098 585898 483334
rect 585342 443418 585578 443654
rect 585662 443418 585898 443654
rect 585342 443098 585578 443334
rect 585662 443098 585898 443334
rect 585342 403418 585578 403654
rect 585662 403418 585898 403654
rect 585342 403098 585578 403334
rect 585662 403098 585898 403334
rect 585342 363418 585578 363654
rect 585662 363418 585898 363654
rect 585342 363098 585578 363334
rect 585662 363098 585898 363334
rect 585342 323418 585578 323654
rect 585662 323418 585898 323654
rect 585342 323098 585578 323334
rect 585662 323098 585898 323334
rect 585342 283418 585578 283654
rect 585662 283418 585898 283654
rect 585342 283098 585578 283334
rect 585662 283098 585898 283334
rect 585342 243418 585578 243654
rect 585662 243418 585898 243654
rect 585342 243098 585578 243334
rect 585662 243098 585898 243334
rect 585342 203418 585578 203654
rect 585662 203418 585898 203654
rect 585342 203098 585578 203334
rect 585662 203098 585898 203334
rect 585342 163418 585578 163654
rect 585662 163418 585898 163654
rect 585342 163098 585578 163334
rect 585662 163098 585898 163334
rect 585342 123418 585578 123654
rect 585662 123418 585898 123654
rect 585342 123098 585578 123334
rect 585662 123098 585898 123334
rect 585342 83418 585578 83654
rect 585662 83418 585898 83654
rect 585342 83098 585578 83334
rect 585662 83098 585898 83334
rect 585342 43418 585578 43654
rect 585662 43418 585898 43654
rect 585342 43098 585578 43334
rect 585662 43098 585898 43334
rect 585342 3418 585578 3654
rect 585662 3418 585898 3654
rect 585342 3098 585578 3334
rect 585662 3098 585898 3334
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 588452 687138 588688 687374
rect 588772 687138 589008 687374
rect 588452 686818 588688 687054
rect 588772 686818 589008 687054
rect 588452 647138 588688 647374
rect 588772 647138 589008 647374
rect 588452 646818 588688 647054
rect 588772 646818 589008 647054
rect 588452 607138 588688 607374
rect 588772 607138 589008 607374
rect 588452 606818 588688 607054
rect 588772 606818 589008 607054
rect 588452 567138 588688 567374
rect 588772 567138 589008 567374
rect 588452 566818 588688 567054
rect 588772 566818 589008 567054
rect 588452 527138 588688 527374
rect 588772 527138 589008 527374
rect 588452 526818 588688 527054
rect 588772 526818 589008 527054
rect 588452 487138 588688 487374
rect 588772 487138 589008 487374
rect 588452 486818 588688 487054
rect 588772 486818 589008 487054
rect 588452 447138 588688 447374
rect 588772 447138 589008 447374
rect 588452 446818 588688 447054
rect 588772 446818 589008 447054
rect 588452 407138 588688 407374
rect 588772 407138 589008 407374
rect 588452 406818 588688 407054
rect 588772 406818 589008 407054
rect 588452 367138 588688 367374
rect 588772 367138 589008 367374
rect 588452 366818 588688 367054
rect 588772 366818 589008 367054
rect 588452 327138 588688 327374
rect 588772 327138 589008 327374
rect 588452 326818 588688 327054
rect 588772 326818 589008 327054
rect 588452 287138 588688 287374
rect 588772 287138 589008 287374
rect 588452 286818 588688 287054
rect 588772 286818 589008 287054
rect 588452 247138 588688 247374
rect 588772 247138 589008 247374
rect 588452 246818 588688 247054
rect 588772 246818 589008 247054
rect 588452 207138 588688 207374
rect 588772 207138 589008 207374
rect 588452 206818 588688 207054
rect 588772 206818 589008 207054
rect 588452 167138 588688 167374
rect 588772 167138 589008 167374
rect 588452 166818 588688 167054
rect 588772 166818 589008 167054
rect 588452 127138 588688 127374
rect 588772 127138 589008 127374
rect 588452 126818 588688 127054
rect 588772 126818 589008 127054
rect 588452 87138 588688 87374
rect 588772 87138 589008 87374
rect 588452 86818 588688 87054
rect 588772 86818 589008 87054
rect 588452 47138 588688 47374
rect 588772 47138 589008 47374
rect 588452 46818 588688 47054
rect 588772 46818 589008 47054
rect 588452 7138 588688 7374
rect 588772 7138 589008 7374
rect 588452 6818 588688 7054
rect 588772 6818 589008 7054
rect 588452 -3692 588688 -3456
rect 588772 -3692 589008 -3456
rect 588452 -4012 588688 -3776
rect 588772 -4012 589008 -3776
rect 591562 690858 591798 691094
rect 591882 690858 592118 691094
rect 591562 690538 591798 690774
rect 591882 690538 592118 690774
rect 591562 650858 591798 651094
rect 591882 650858 592118 651094
rect 591562 650538 591798 650774
rect 591882 650538 592118 650774
rect 591562 610858 591798 611094
rect 591882 610858 592118 611094
rect 591562 610538 591798 610774
rect 591882 610538 592118 610774
rect 591562 570858 591798 571094
rect 591882 570858 592118 571094
rect 591562 570538 591798 570774
rect 591882 570538 592118 570774
rect 591562 530858 591798 531094
rect 591882 530858 592118 531094
rect 591562 530538 591798 530774
rect 591882 530538 592118 530774
rect 591562 490858 591798 491094
rect 591882 490858 592118 491094
rect 591562 490538 591798 490774
rect 591882 490538 592118 490774
rect 591562 450858 591798 451094
rect 591882 450858 592118 451094
rect 591562 450538 591798 450774
rect 591882 450538 592118 450774
rect 591562 410858 591798 411094
rect 591882 410858 592118 411094
rect 591562 410538 591798 410774
rect 591882 410538 592118 410774
rect 591562 370858 591798 371094
rect 591882 370858 592118 371094
rect 591562 370538 591798 370774
rect 591882 370538 592118 370774
rect 591562 330858 591798 331094
rect 591882 330858 592118 331094
rect 591562 330538 591798 330774
rect 591882 330538 592118 330774
rect 591562 290858 591798 291094
rect 591882 290858 592118 291094
rect 591562 290538 591798 290774
rect 591882 290538 592118 290774
rect 591562 250858 591798 251094
rect 591882 250858 592118 251094
rect 591562 250538 591798 250774
rect 591882 250538 592118 250774
rect 591562 210858 591798 211094
rect 591882 210858 592118 211094
rect 591562 210538 591798 210774
rect 591882 210538 592118 210774
rect 591562 170858 591798 171094
rect 591882 170858 592118 171094
rect 591562 170538 591798 170774
rect 591882 170538 592118 170774
rect 591562 130858 591798 131094
rect 591882 130858 592118 131094
rect 591562 130538 591798 130774
rect 591882 130538 592118 130774
rect 591562 90858 591798 91094
rect 591882 90858 592118 91094
rect 591562 90538 591798 90774
rect 591882 90538 592118 90774
rect 591562 50858 591798 51094
rect 591882 50858 592118 51094
rect 591562 50538 591798 50774
rect 591882 50538 592118 50774
rect 591562 10858 591798 11094
rect 591882 10858 592118 11094
rect 591562 10538 591798 10774
rect 591882 10538 592118 10774
rect 591562 -6802 591798 -6566
rect 591882 -6802 592118 -6566
rect 591562 -7122 591798 -6886
rect 591882 -7122 592118 -6886
rect 594672 694578 594908 694814
rect 594992 694578 595228 694814
rect 594672 694258 594908 694494
rect 594992 694258 595228 694494
rect 594672 654578 594908 654814
rect 594992 654578 595228 654814
rect 594672 654258 594908 654494
rect 594992 654258 595228 654494
rect 594672 614578 594908 614814
rect 594992 614578 595228 614814
rect 594672 614258 594908 614494
rect 594992 614258 595228 614494
rect 594672 574578 594908 574814
rect 594992 574578 595228 574814
rect 594672 574258 594908 574494
rect 594992 574258 595228 574494
rect 594672 534578 594908 534814
rect 594992 534578 595228 534814
rect 594672 534258 594908 534494
rect 594992 534258 595228 534494
rect 594672 494578 594908 494814
rect 594992 494578 595228 494814
rect 594672 494258 594908 494494
rect 594992 494258 595228 494494
rect 594672 454578 594908 454814
rect 594992 454578 595228 454814
rect 594672 454258 594908 454494
rect 594992 454258 595228 454494
rect 594672 414578 594908 414814
rect 594992 414578 595228 414814
rect 594672 414258 594908 414494
rect 594992 414258 595228 414494
rect 594672 374578 594908 374814
rect 594992 374578 595228 374814
rect 594672 374258 594908 374494
rect 594992 374258 595228 374494
rect 594672 334578 594908 334814
rect 594992 334578 595228 334814
rect 594672 334258 594908 334494
rect 594992 334258 595228 334494
rect 594672 294578 594908 294814
rect 594992 294578 595228 294814
rect 594672 294258 594908 294494
rect 594992 294258 595228 294494
rect 594672 254578 594908 254814
rect 594992 254578 595228 254814
rect 594672 254258 594908 254494
rect 594992 254258 595228 254494
rect 594672 214578 594908 214814
rect 594992 214578 595228 214814
rect 594672 214258 594908 214494
rect 594992 214258 595228 214494
rect 594672 174578 594908 174814
rect 594992 174578 595228 174814
rect 594672 174258 594908 174494
rect 594992 174258 595228 174494
rect 594672 134578 594908 134814
rect 594992 134578 595228 134814
rect 594672 134258 594908 134494
rect 594992 134258 595228 134494
rect 594672 94578 594908 94814
rect 594992 94578 595228 94814
rect 594672 94258 594908 94494
rect 594992 94258 595228 94494
rect 594672 54578 594908 54814
rect 594992 54578 595228 54814
rect 594672 54258 594908 54494
rect 594992 54258 595228 54494
rect 594672 14578 594908 14814
rect 594992 14578 595228 14814
rect 594672 14258 594908 14494
rect 594992 14258 595228 14494
rect 594672 -9912 594908 -9676
rect 594992 -9912 595228 -9676
rect 594672 -10232 594908 -9996
rect 594992 -10232 595228 -9996
rect 597782 698298 598018 698534
rect 598102 698298 598338 698534
rect 597782 697978 598018 698214
rect 598102 697978 598338 698214
rect 597782 658298 598018 658534
rect 598102 658298 598338 658534
rect 597782 657978 598018 658214
rect 598102 657978 598338 658214
rect 597782 618298 598018 618534
rect 598102 618298 598338 618534
rect 597782 617978 598018 618214
rect 598102 617978 598338 618214
rect 597782 578298 598018 578534
rect 598102 578298 598338 578534
rect 597782 577978 598018 578214
rect 598102 577978 598338 578214
rect 597782 538298 598018 538534
rect 598102 538298 598338 538534
rect 597782 537978 598018 538214
rect 598102 537978 598338 538214
rect 597782 498298 598018 498534
rect 598102 498298 598338 498534
rect 597782 497978 598018 498214
rect 598102 497978 598338 498214
rect 597782 458298 598018 458534
rect 598102 458298 598338 458534
rect 597782 457978 598018 458214
rect 598102 457978 598338 458214
rect 597782 418298 598018 418534
rect 598102 418298 598338 418534
rect 597782 417978 598018 418214
rect 598102 417978 598338 418214
rect 597782 378298 598018 378534
rect 598102 378298 598338 378534
rect 597782 377978 598018 378214
rect 598102 377978 598338 378214
rect 597782 338298 598018 338534
rect 598102 338298 598338 338534
rect 597782 337978 598018 338214
rect 598102 337978 598338 338214
rect 597782 298298 598018 298534
rect 598102 298298 598338 298534
rect 597782 297978 598018 298214
rect 598102 297978 598338 298214
rect 597782 258298 598018 258534
rect 598102 258298 598338 258534
rect 597782 257978 598018 258214
rect 598102 257978 598338 258214
rect 597782 218298 598018 218534
rect 598102 218298 598338 218534
rect 597782 217978 598018 218214
rect 598102 217978 598338 218214
rect 597782 178298 598018 178534
rect 598102 178298 598338 178534
rect 597782 177978 598018 178214
rect 598102 177978 598338 178214
rect 597782 138298 598018 138534
rect 598102 138298 598338 138534
rect 597782 137978 598018 138214
rect 598102 137978 598338 138214
rect 597782 98298 598018 98534
rect 598102 98298 598338 98534
rect 597782 97978 598018 98214
rect 598102 97978 598338 98214
rect 597782 58298 598018 58534
rect 598102 58298 598338 58534
rect 597782 57978 598018 58214
rect 598102 57978 598338 58214
rect 597782 18298 598018 18534
rect 598102 18298 598338 18534
rect 597782 17978 598018 18214
rect 598102 17978 598338 18214
rect 597782 -13022 598018 -12786
rect 598102 -13022 598338 -12786
rect 597782 -13342 598018 -13106
rect 598102 -13342 598338 -13106
rect 600892 662018 601128 662254
rect 601212 662018 601448 662254
rect 600892 661698 601128 661934
rect 601212 661698 601448 661934
rect 600892 622018 601128 622254
rect 601212 622018 601448 622254
rect 600892 621698 601128 621934
rect 601212 621698 601448 621934
rect 600892 582018 601128 582254
rect 601212 582018 601448 582254
rect 600892 581698 601128 581934
rect 601212 581698 601448 581934
rect 600892 542018 601128 542254
rect 601212 542018 601448 542254
rect 600892 541698 601128 541934
rect 601212 541698 601448 541934
rect 600892 502018 601128 502254
rect 601212 502018 601448 502254
rect 600892 501698 601128 501934
rect 601212 501698 601448 501934
rect 600892 462018 601128 462254
rect 601212 462018 601448 462254
rect 600892 461698 601128 461934
rect 601212 461698 601448 461934
rect 600892 422018 601128 422254
rect 601212 422018 601448 422254
rect 600892 421698 601128 421934
rect 601212 421698 601448 421934
rect 600892 382018 601128 382254
rect 601212 382018 601448 382254
rect 600892 381698 601128 381934
rect 601212 381698 601448 381934
rect 600892 342018 601128 342254
rect 601212 342018 601448 342254
rect 600892 341698 601128 341934
rect 601212 341698 601448 341934
rect 600892 302018 601128 302254
rect 601212 302018 601448 302254
rect 600892 301698 601128 301934
rect 601212 301698 601448 301934
rect 600892 262018 601128 262254
rect 601212 262018 601448 262254
rect 600892 261698 601128 261934
rect 601212 261698 601448 261934
rect 600892 222018 601128 222254
rect 601212 222018 601448 222254
rect 600892 221698 601128 221934
rect 601212 221698 601448 221934
rect 600892 182018 601128 182254
rect 601212 182018 601448 182254
rect 600892 181698 601128 181934
rect 601212 181698 601448 181934
rect 600892 142018 601128 142254
rect 601212 142018 601448 142254
rect 600892 141698 601128 141934
rect 601212 141698 601448 141934
rect 600892 102018 601128 102254
rect 601212 102018 601448 102254
rect 600892 101698 601128 101934
rect 601212 101698 601448 101934
rect 600892 62018 601128 62254
rect 601212 62018 601448 62254
rect 600892 61698 601128 61934
rect 601212 61698 601448 61934
rect 600892 22018 601128 22254
rect 601212 22018 601448 22254
rect 600892 21698 601128 21934
rect 601212 21698 601448 21934
rect 580626 -16132 580862 -15896
rect 580946 -16132 581182 -15896
rect 580626 -16452 580862 -16216
rect 580946 -16452 581182 -16216
rect -20634 -19242 -20398 -19006
rect -20314 -19242 -20078 -19006
rect -20634 -19562 -20398 -19326
rect -20314 -19562 -20078 -19326
rect -23744 -22352 -23508 -22116
rect -23424 -22352 -23188 -22116
rect -23744 -22672 -23508 -22436
rect -23424 -22672 -23188 -22436
rect 600892 -16132 601128 -15896
rect 601212 -16132 601448 -15896
rect 600892 -16452 601128 -16216
rect 601212 -16452 601448 -16216
rect 604002 665738 604238 665974
rect 604322 665738 604558 665974
rect 604002 665418 604238 665654
rect 604322 665418 604558 665654
rect 604002 625738 604238 625974
rect 604322 625738 604558 625974
rect 604002 625418 604238 625654
rect 604322 625418 604558 625654
rect 604002 585738 604238 585974
rect 604322 585738 604558 585974
rect 604002 585418 604238 585654
rect 604322 585418 604558 585654
rect 604002 545738 604238 545974
rect 604322 545738 604558 545974
rect 604002 545418 604238 545654
rect 604322 545418 604558 545654
rect 604002 505738 604238 505974
rect 604322 505738 604558 505974
rect 604002 505418 604238 505654
rect 604322 505418 604558 505654
rect 604002 465738 604238 465974
rect 604322 465738 604558 465974
rect 604002 465418 604238 465654
rect 604322 465418 604558 465654
rect 604002 425738 604238 425974
rect 604322 425738 604558 425974
rect 604002 425418 604238 425654
rect 604322 425418 604558 425654
rect 604002 385738 604238 385974
rect 604322 385738 604558 385974
rect 604002 385418 604238 385654
rect 604322 385418 604558 385654
rect 604002 345738 604238 345974
rect 604322 345738 604558 345974
rect 604002 345418 604238 345654
rect 604322 345418 604558 345654
rect 604002 305738 604238 305974
rect 604322 305738 604558 305974
rect 604002 305418 604238 305654
rect 604322 305418 604558 305654
rect 604002 265738 604238 265974
rect 604322 265738 604558 265974
rect 604002 265418 604238 265654
rect 604322 265418 604558 265654
rect 604002 225738 604238 225974
rect 604322 225738 604558 225974
rect 604002 225418 604238 225654
rect 604322 225418 604558 225654
rect 604002 185738 604238 185974
rect 604322 185738 604558 185974
rect 604002 185418 604238 185654
rect 604322 185418 604558 185654
rect 604002 145738 604238 145974
rect 604322 145738 604558 145974
rect 604002 145418 604238 145654
rect 604322 145418 604558 145654
rect 604002 105738 604238 105974
rect 604322 105738 604558 105974
rect 604002 105418 604238 105654
rect 604322 105418 604558 105654
rect 604002 65738 604238 65974
rect 604322 65738 604558 65974
rect 604002 65418 604238 65654
rect 604322 65418 604558 65654
rect 604002 25738 604238 25974
rect 604322 25738 604558 25974
rect 604002 25418 604238 25654
rect 604322 25418 604558 25654
rect 604002 -19242 604238 -19006
rect 604322 -19242 604558 -19006
rect 604002 -19562 604238 -19326
rect 604322 -19562 604558 -19326
rect 607112 669458 607348 669694
rect 607432 669458 607668 669694
rect 607112 669138 607348 669374
rect 607432 669138 607668 669374
rect 607112 629458 607348 629694
rect 607432 629458 607668 629694
rect 607112 629138 607348 629374
rect 607432 629138 607668 629374
rect 607112 589458 607348 589694
rect 607432 589458 607668 589694
rect 607112 589138 607348 589374
rect 607432 589138 607668 589374
rect 607112 549458 607348 549694
rect 607432 549458 607668 549694
rect 607112 549138 607348 549374
rect 607432 549138 607668 549374
rect 607112 509458 607348 509694
rect 607432 509458 607668 509694
rect 607112 509138 607348 509374
rect 607432 509138 607668 509374
rect 607112 469458 607348 469694
rect 607432 469458 607668 469694
rect 607112 469138 607348 469374
rect 607432 469138 607668 469374
rect 607112 429458 607348 429694
rect 607432 429458 607668 429694
rect 607112 429138 607348 429374
rect 607432 429138 607668 429374
rect 607112 389458 607348 389694
rect 607432 389458 607668 389694
rect 607112 389138 607348 389374
rect 607432 389138 607668 389374
rect 607112 349458 607348 349694
rect 607432 349458 607668 349694
rect 607112 349138 607348 349374
rect 607432 349138 607668 349374
rect 607112 309458 607348 309694
rect 607432 309458 607668 309694
rect 607112 309138 607348 309374
rect 607432 309138 607668 309374
rect 607112 269458 607348 269694
rect 607432 269458 607668 269694
rect 607112 269138 607348 269374
rect 607432 269138 607668 269374
rect 607112 229458 607348 229694
rect 607432 229458 607668 229694
rect 607112 229138 607348 229374
rect 607432 229138 607668 229374
rect 607112 189458 607348 189694
rect 607432 189458 607668 189694
rect 607112 189138 607348 189374
rect 607432 189138 607668 189374
rect 607112 149458 607348 149694
rect 607432 149458 607668 149694
rect 607112 149138 607348 149374
rect 607432 149138 607668 149374
rect 607112 109458 607348 109694
rect 607432 109458 607668 109694
rect 607112 109138 607348 109374
rect 607432 109138 607668 109374
rect 607112 69458 607348 69694
rect 607432 69458 607668 69694
rect 607112 69138 607348 69374
rect 607432 69138 607668 69374
rect 607112 29458 607348 29694
rect 607432 29458 607668 29694
rect 607112 29138 607348 29374
rect 607432 29138 607668 29374
rect 607112 -22352 607348 -22116
rect 607432 -22352 607668 -22116
rect 607112 -22672 607348 -22436
rect 607432 -22672 607668 -22436
<< metal5 >>
rect -23776 726608 607700 726640
rect -23776 726372 -23744 726608
rect -23508 726372 -23424 726608
rect -23188 726372 607112 726608
rect 607348 726372 607432 726608
rect 607668 726372 607700 726608
rect -23776 726288 607700 726372
rect -23776 726052 -23744 726288
rect -23508 726052 -23424 726288
rect -23188 726052 607112 726288
rect 607348 726052 607432 726288
rect 607668 726052 607700 726288
rect -23776 726020 607700 726052
rect -20666 723498 604590 723530
rect -20666 723262 -20634 723498
rect -20398 723262 -20314 723498
rect -20078 723262 604002 723498
rect 604238 723262 604322 723498
rect 604558 723262 604590 723498
rect -20666 723178 604590 723262
rect -20666 722942 -20634 723178
rect -20398 722942 -20314 723178
rect -20078 722942 604002 723178
rect 604238 722942 604322 723178
rect 604558 722942 604590 723178
rect -20666 722910 604590 722942
rect -17556 720388 601480 720420
rect -17556 720152 -17524 720388
rect -17288 720152 -17204 720388
rect -16968 720152 580626 720388
rect 580862 720152 580946 720388
rect 581182 720152 600892 720388
rect 601128 720152 601212 720388
rect 601448 720152 601480 720388
rect -17556 720068 601480 720152
rect -17556 719832 -17524 720068
rect -17288 719832 -17204 720068
rect -16968 719832 580626 720068
rect 580862 719832 580946 720068
rect 581182 719832 600892 720068
rect 601128 719832 601212 720068
rect 601448 719832 601480 720068
rect -17556 719800 601480 719832
rect -14446 717278 598370 717310
rect -14446 717042 -14414 717278
rect -14178 717042 -14094 717278
rect -13858 717042 597782 717278
rect 598018 717042 598102 717278
rect 598338 717042 598370 717278
rect -14446 716958 598370 717042
rect -14446 716722 -14414 716958
rect -14178 716722 -14094 716958
rect -13858 716722 597782 716958
rect 598018 716722 598102 716958
rect 598338 716722 598370 716958
rect -14446 716690 598370 716722
rect -11336 714168 595260 714200
rect -11336 713932 -11304 714168
rect -11068 713932 -10984 714168
rect -10748 713932 594672 714168
rect 594908 713932 594992 714168
rect 595228 713932 595260 714168
rect -11336 713848 595260 713932
rect -11336 713612 -11304 713848
rect -11068 713612 -10984 713848
rect -10748 713612 594672 713848
rect 594908 713612 594992 713848
rect 595228 713612 595260 713848
rect -11336 713580 595260 713612
rect -8226 711058 592150 711090
rect -8226 710822 -8194 711058
rect -7958 710822 -7874 711058
rect -7638 710822 591562 711058
rect 591798 710822 591882 711058
rect 592118 710822 592150 711058
rect -8226 710738 592150 710822
rect -8226 710502 -8194 710738
rect -7958 710502 -7874 710738
rect -7638 710502 591562 710738
rect 591798 710502 591882 710738
rect 592118 710502 592150 710738
rect -8226 710470 592150 710502
rect -5116 707948 589040 707980
rect -5116 707712 -5084 707948
rect -4848 707712 -4764 707948
rect -4528 707712 588452 707948
rect 588688 707712 588772 707948
rect 589008 707712 589040 707948
rect -5116 707628 589040 707712
rect -5116 707392 -5084 707628
rect -4848 707392 -4764 707628
rect -4528 707392 588452 707628
rect 588688 707392 588772 707628
rect 589008 707392 589040 707628
rect -5116 707360 589040 707392
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -23776 698534 607700 698566
rect -23776 698298 -14414 698534
rect -14178 698298 -14094 698534
rect -13858 698298 597782 698534
rect 598018 698298 598102 698534
rect 598338 698298 607700 698534
rect -23776 698214 607700 698298
rect -23776 697978 -14414 698214
rect -14178 697978 -14094 698214
rect -13858 697978 597782 698214
rect 598018 697978 598102 698214
rect 598338 697978 607700 698214
rect -23776 697946 607700 697978
rect -23776 694814 607700 694846
rect -23776 694578 -11304 694814
rect -11068 694578 -10984 694814
rect -10748 694578 594672 694814
rect 594908 694578 594992 694814
rect 595228 694578 607700 694814
rect -23776 694494 607700 694578
rect -23776 694258 -11304 694494
rect -11068 694258 -10984 694494
rect -10748 694258 594672 694494
rect 594908 694258 594992 694494
rect 595228 694258 607700 694494
rect -23776 694226 607700 694258
rect 7852 693716 8456 693748
rect 7852 693480 7876 693716
rect 8112 693480 8196 693716
rect 8432 693480 8456 693716
rect 7852 693396 8456 693480
rect 7852 693160 7876 693396
rect 8112 693160 8196 693396
rect 8432 693160 8456 693396
rect 7852 693128 8456 693160
rect 38008 693716 38612 693748
rect 38008 693480 38032 693716
rect 38268 693480 38352 693716
rect 38588 693480 38612 693716
rect 38008 693396 38612 693480
rect 38008 693160 38032 693396
rect 38268 693160 38352 693396
rect 38588 693160 38612 693396
rect 38008 693128 38612 693160
rect 74008 693716 74612 693748
rect 74008 693480 74032 693716
rect 74268 693480 74352 693716
rect 74588 693480 74612 693716
rect 74008 693396 74612 693480
rect 74008 693160 74032 693396
rect 74268 693160 74352 693396
rect 74588 693160 74612 693396
rect 74008 693128 74612 693160
rect 110008 693716 110612 693748
rect 110008 693480 110032 693716
rect 110268 693480 110352 693716
rect 110588 693480 110612 693716
rect 110008 693396 110612 693480
rect 110008 693160 110032 693396
rect 110268 693160 110352 693396
rect 110588 693160 110612 693396
rect 110008 693128 110612 693160
rect 146008 693716 146612 693748
rect 146008 693480 146032 693716
rect 146268 693480 146352 693716
rect 146588 693480 146612 693716
rect 146008 693396 146612 693480
rect 146008 693160 146032 693396
rect 146268 693160 146352 693396
rect 146588 693160 146612 693396
rect 146008 693128 146612 693160
rect 182008 693716 182612 693748
rect 182008 693480 182032 693716
rect 182268 693480 182352 693716
rect 182588 693480 182612 693716
rect 182008 693396 182612 693480
rect 182008 693160 182032 693396
rect 182268 693160 182352 693396
rect 182588 693160 182612 693396
rect 182008 693128 182612 693160
rect 218008 693716 218612 693748
rect 218008 693480 218032 693716
rect 218268 693480 218352 693716
rect 218588 693480 218612 693716
rect 218008 693396 218612 693480
rect 218008 693160 218032 693396
rect 218268 693160 218352 693396
rect 218588 693160 218612 693396
rect 218008 693128 218612 693160
rect 254008 693716 254612 693748
rect 254008 693480 254032 693716
rect 254268 693480 254352 693716
rect 254588 693480 254612 693716
rect 254008 693396 254612 693480
rect 254008 693160 254032 693396
rect 254268 693160 254352 693396
rect 254588 693160 254612 693396
rect 254008 693128 254612 693160
rect 290008 693716 290612 693748
rect 290008 693480 290032 693716
rect 290268 693480 290352 693716
rect 290588 693480 290612 693716
rect 290008 693396 290612 693480
rect 290008 693160 290032 693396
rect 290268 693160 290352 693396
rect 290588 693160 290612 693396
rect 290008 693128 290612 693160
rect 326008 693716 326612 693748
rect 326008 693480 326032 693716
rect 326268 693480 326352 693716
rect 326588 693480 326612 693716
rect 326008 693396 326612 693480
rect 326008 693160 326032 693396
rect 326268 693160 326352 693396
rect 326588 693160 326612 693396
rect 326008 693128 326612 693160
rect 362008 693716 362612 693748
rect 362008 693480 362032 693716
rect 362268 693480 362352 693716
rect 362588 693480 362612 693716
rect 362008 693396 362612 693480
rect 362008 693160 362032 693396
rect 362268 693160 362352 693396
rect 362588 693160 362612 693396
rect 362008 693128 362612 693160
rect 398008 693716 398612 693748
rect 398008 693480 398032 693716
rect 398268 693480 398352 693716
rect 398588 693480 398612 693716
rect 398008 693396 398612 693480
rect 398008 693160 398032 693396
rect 398268 693160 398352 693396
rect 398588 693160 398612 693396
rect 398008 693128 398612 693160
rect 434008 693716 434612 693748
rect 434008 693480 434032 693716
rect 434268 693480 434352 693716
rect 434588 693480 434612 693716
rect 434008 693396 434612 693480
rect 434008 693160 434032 693396
rect 434268 693160 434352 693396
rect 434588 693160 434612 693396
rect 434008 693128 434612 693160
rect 470008 693716 470612 693748
rect 470008 693480 470032 693716
rect 470268 693480 470352 693716
rect 470588 693480 470612 693716
rect 470008 693396 470612 693480
rect 470008 693160 470032 693396
rect 470268 693160 470352 693396
rect 470588 693160 470612 693396
rect 470008 693128 470612 693160
rect 506008 693716 506612 693748
rect 506008 693480 506032 693716
rect 506268 693480 506352 693716
rect 506588 693480 506612 693716
rect 506008 693396 506612 693480
rect 506008 693160 506032 693396
rect 506268 693160 506352 693396
rect 506588 693160 506612 693396
rect 506008 693128 506612 693160
rect 542008 693716 542612 693748
rect 542008 693480 542032 693716
rect 542268 693480 542352 693716
rect 542588 693480 542612 693716
rect 542008 693396 542612 693480
rect 542008 693160 542032 693396
rect 542268 693160 542352 693396
rect 542588 693160 542612 693396
rect 542008 693128 542612 693160
rect 571508 693716 572112 693748
rect 571508 693480 571532 693716
rect 571768 693480 571852 693716
rect 572088 693480 572112 693716
rect 571508 693396 572112 693480
rect 571508 693160 571532 693396
rect 571768 693160 571852 693396
rect 572088 693160 572112 693396
rect 571508 693128 572112 693160
rect 9092 692476 9696 692508
rect 9092 692240 9116 692476
rect 9352 692240 9436 692476
rect 9672 692240 9696 692476
rect 9092 692156 9696 692240
rect 9092 691920 9116 692156
rect 9352 691920 9436 692156
rect 9672 691920 9696 692156
rect 9092 691888 9696 691920
rect 56628 692476 57232 692508
rect 56628 692240 56652 692476
rect 56888 692240 56972 692476
rect 57208 692240 57232 692476
rect 56628 692156 57232 692240
rect 56628 691920 56652 692156
rect 56888 691920 56972 692156
rect 57208 691920 57232 692156
rect 56628 691888 57232 691920
rect 92628 692476 93232 692508
rect 92628 692240 92652 692476
rect 92888 692240 92972 692476
rect 93208 692240 93232 692476
rect 92628 692156 93232 692240
rect 92628 691920 92652 692156
rect 92888 691920 92972 692156
rect 93208 691920 93232 692156
rect 92628 691888 93232 691920
rect 128628 692476 129232 692508
rect 128628 692240 128652 692476
rect 128888 692240 128972 692476
rect 129208 692240 129232 692476
rect 128628 692156 129232 692240
rect 128628 691920 128652 692156
rect 128888 691920 128972 692156
rect 129208 691920 129232 692156
rect 128628 691888 129232 691920
rect 164628 692476 165232 692508
rect 164628 692240 164652 692476
rect 164888 692240 164972 692476
rect 165208 692240 165232 692476
rect 164628 692156 165232 692240
rect 164628 691920 164652 692156
rect 164888 691920 164972 692156
rect 165208 691920 165232 692156
rect 164628 691888 165232 691920
rect 200628 692476 201232 692508
rect 200628 692240 200652 692476
rect 200888 692240 200972 692476
rect 201208 692240 201232 692476
rect 200628 692156 201232 692240
rect 200628 691920 200652 692156
rect 200888 691920 200972 692156
rect 201208 691920 201232 692156
rect 200628 691888 201232 691920
rect 236628 692476 237232 692508
rect 236628 692240 236652 692476
rect 236888 692240 236972 692476
rect 237208 692240 237232 692476
rect 236628 692156 237232 692240
rect 236628 691920 236652 692156
rect 236888 691920 236972 692156
rect 237208 691920 237232 692156
rect 236628 691888 237232 691920
rect 272628 692476 273232 692508
rect 272628 692240 272652 692476
rect 272888 692240 272972 692476
rect 273208 692240 273232 692476
rect 272628 692156 273232 692240
rect 272628 691920 272652 692156
rect 272888 691920 272972 692156
rect 273208 691920 273232 692156
rect 272628 691888 273232 691920
rect 308628 692476 309232 692508
rect 308628 692240 308652 692476
rect 308888 692240 308972 692476
rect 309208 692240 309232 692476
rect 308628 692156 309232 692240
rect 308628 691920 308652 692156
rect 308888 691920 308972 692156
rect 309208 691920 309232 692156
rect 308628 691888 309232 691920
rect 344628 692476 345232 692508
rect 344628 692240 344652 692476
rect 344888 692240 344972 692476
rect 345208 692240 345232 692476
rect 344628 692156 345232 692240
rect 344628 691920 344652 692156
rect 344888 691920 344972 692156
rect 345208 691920 345232 692156
rect 344628 691888 345232 691920
rect 380628 692476 381232 692508
rect 380628 692240 380652 692476
rect 380888 692240 380972 692476
rect 381208 692240 381232 692476
rect 380628 692156 381232 692240
rect 380628 691920 380652 692156
rect 380888 691920 380972 692156
rect 381208 691920 381232 692156
rect 380628 691888 381232 691920
rect 416628 692476 417232 692508
rect 416628 692240 416652 692476
rect 416888 692240 416972 692476
rect 417208 692240 417232 692476
rect 416628 692156 417232 692240
rect 416628 691920 416652 692156
rect 416888 691920 416972 692156
rect 417208 691920 417232 692156
rect 416628 691888 417232 691920
rect 452628 692476 453232 692508
rect 452628 692240 452652 692476
rect 452888 692240 452972 692476
rect 453208 692240 453232 692476
rect 452628 692156 453232 692240
rect 452628 691920 452652 692156
rect 452888 691920 452972 692156
rect 453208 691920 453232 692156
rect 452628 691888 453232 691920
rect 488628 692476 489232 692508
rect 488628 692240 488652 692476
rect 488888 692240 488972 692476
rect 489208 692240 489232 692476
rect 488628 692156 489232 692240
rect 488628 691920 488652 692156
rect 488888 691920 488972 692156
rect 489208 691920 489232 692156
rect 488628 691888 489232 691920
rect 524628 692476 525232 692508
rect 524628 692240 524652 692476
rect 524888 692240 524972 692476
rect 525208 692240 525232 692476
rect 524628 692156 525232 692240
rect 524628 691920 524652 692156
rect 524888 691920 524972 692156
rect 525208 691920 525232 692156
rect 524628 691888 525232 691920
rect 560628 692476 561232 692508
rect 560628 692240 560652 692476
rect 560888 692240 560972 692476
rect 561208 692240 561232 692476
rect 560628 692156 561232 692240
rect 560628 691920 560652 692156
rect 560888 691920 560972 692156
rect 561208 691920 561232 692156
rect 560628 691888 561232 691920
rect 570268 692476 570872 692508
rect 570268 692240 570292 692476
rect 570528 692240 570612 692476
rect 570848 692240 570872 692476
rect 570268 692156 570872 692240
rect 570268 691920 570292 692156
rect 570528 691920 570612 692156
rect 570848 691920 570872 692156
rect 570268 691888 570872 691920
rect -23776 691094 607700 691126
rect -23776 690858 -8194 691094
rect -7958 690858 -7874 691094
rect -7638 690858 591562 691094
rect 591798 690858 591882 691094
rect 592118 690858 607700 691094
rect -23776 690774 607700 690858
rect -23776 690538 -8194 690774
rect -7958 690538 -7874 690774
rect -7638 690538 591562 690774
rect 591798 690538 591882 690774
rect 592118 690538 607700 690774
rect -23776 690506 607700 690538
rect -23776 687374 607700 687406
rect -23776 687138 -5084 687374
rect -4848 687138 -4764 687374
rect -4528 687138 7876 687374
rect 8112 687138 8196 687374
rect 8432 687138 38032 687374
rect 38268 687138 38352 687374
rect 38588 687138 74032 687374
rect 74268 687138 74352 687374
rect 74588 687138 110032 687374
rect 110268 687138 110352 687374
rect 110588 687138 146032 687374
rect 146268 687138 146352 687374
rect 146588 687138 182032 687374
rect 182268 687138 182352 687374
rect 182588 687138 218032 687374
rect 218268 687138 218352 687374
rect 218588 687138 254032 687374
rect 254268 687138 254352 687374
rect 254588 687138 290032 687374
rect 290268 687138 290352 687374
rect 290588 687138 326032 687374
rect 326268 687138 326352 687374
rect 326588 687138 362032 687374
rect 362268 687138 362352 687374
rect 362588 687138 398032 687374
rect 398268 687138 398352 687374
rect 398588 687138 434032 687374
rect 434268 687138 434352 687374
rect 434588 687138 470032 687374
rect 470268 687138 470352 687374
rect 470588 687138 506032 687374
rect 506268 687138 506352 687374
rect 506588 687138 542032 687374
rect 542268 687138 542352 687374
rect 542588 687138 571532 687374
rect 571768 687138 571852 687374
rect 572088 687138 588452 687374
rect 588688 687138 588772 687374
rect 589008 687138 607700 687374
rect -23776 687054 607700 687138
rect -23776 686818 -5084 687054
rect -4848 686818 -4764 687054
rect -4528 686818 7876 687054
rect 8112 686818 8196 687054
rect 8432 686818 38032 687054
rect 38268 686818 38352 687054
rect 38588 686818 74032 687054
rect 74268 686818 74352 687054
rect 74588 686818 110032 687054
rect 110268 686818 110352 687054
rect 110588 686818 146032 687054
rect 146268 686818 146352 687054
rect 146588 686818 182032 687054
rect 182268 686818 182352 687054
rect 182588 686818 218032 687054
rect 218268 686818 218352 687054
rect 218588 686818 254032 687054
rect 254268 686818 254352 687054
rect 254588 686818 290032 687054
rect 290268 686818 290352 687054
rect 290588 686818 326032 687054
rect 326268 686818 326352 687054
rect 326588 686818 362032 687054
rect 362268 686818 362352 687054
rect 362588 686818 398032 687054
rect 398268 686818 398352 687054
rect 398588 686818 434032 687054
rect 434268 686818 434352 687054
rect 434588 686818 470032 687054
rect 470268 686818 470352 687054
rect 470588 686818 506032 687054
rect 506268 686818 506352 687054
rect 506588 686818 542032 687054
rect 542268 686818 542352 687054
rect 542588 686818 571532 687054
rect 571768 686818 571852 687054
rect 572088 686818 588452 687054
rect 588688 686818 588772 687054
rect 589008 686818 607700 687054
rect -23776 686786 607700 686818
rect -23776 683654 607700 683686
rect -23776 683418 -1974 683654
rect -1738 683418 -1654 683654
rect -1418 683418 9116 683654
rect 9352 683418 9436 683654
rect 9672 683418 56652 683654
rect 56888 683418 56972 683654
rect 57208 683418 92652 683654
rect 92888 683418 92972 683654
rect 93208 683418 128652 683654
rect 128888 683418 128972 683654
rect 129208 683418 164652 683654
rect 164888 683418 164972 683654
rect 165208 683418 200652 683654
rect 200888 683418 200972 683654
rect 201208 683418 236652 683654
rect 236888 683418 236972 683654
rect 237208 683418 272652 683654
rect 272888 683418 272972 683654
rect 273208 683418 308652 683654
rect 308888 683418 308972 683654
rect 309208 683418 344652 683654
rect 344888 683418 344972 683654
rect 345208 683418 380652 683654
rect 380888 683418 380972 683654
rect 381208 683418 416652 683654
rect 416888 683418 416972 683654
rect 417208 683418 452652 683654
rect 452888 683418 452972 683654
rect 453208 683418 488652 683654
rect 488888 683418 488972 683654
rect 489208 683418 524652 683654
rect 524888 683418 524972 683654
rect 525208 683418 560652 683654
rect 560888 683418 560972 683654
rect 561208 683418 570292 683654
rect 570528 683418 570612 683654
rect 570848 683418 585342 683654
rect 585578 683418 585662 683654
rect 585898 683418 607700 683654
rect -23776 683334 607700 683418
rect -23776 683098 -1974 683334
rect -1738 683098 -1654 683334
rect -1418 683098 9116 683334
rect 9352 683098 9436 683334
rect 9672 683098 56652 683334
rect 56888 683098 56972 683334
rect 57208 683098 92652 683334
rect 92888 683098 92972 683334
rect 93208 683098 128652 683334
rect 128888 683098 128972 683334
rect 129208 683098 164652 683334
rect 164888 683098 164972 683334
rect 165208 683098 200652 683334
rect 200888 683098 200972 683334
rect 201208 683098 236652 683334
rect 236888 683098 236972 683334
rect 237208 683098 272652 683334
rect 272888 683098 272972 683334
rect 273208 683098 308652 683334
rect 308888 683098 308972 683334
rect 309208 683098 344652 683334
rect 344888 683098 344972 683334
rect 345208 683098 380652 683334
rect 380888 683098 380972 683334
rect 381208 683098 416652 683334
rect 416888 683098 416972 683334
rect 417208 683098 452652 683334
rect 452888 683098 452972 683334
rect 453208 683098 488652 683334
rect 488888 683098 488972 683334
rect 489208 683098 524652 683334
rect 524888 683098 524972 683334
rect 525208 683098 560652 683334
rect 560888 683098 560972 683334
rect 561208 683098 570292 683334
rect 570528 683098 570612 683334
rect 570848 683098 585342 683334
rect 585578 683098 585662 683334
rect 585898 683098 607700 683334
rect -23776 683066 607700 683098
rect -23776 669694 607700 669726
rect -23776 669458 -23744 669694
rect -23508 669458 -23424 669694
rect -23188 669458 607112 669694
rect 607348 669458 607432 669694
rect 607668 669458 607700 669694
rect -23776 669374 607700 669458
rect -23776 669138 -23744 669374
rect -23508 669138 -23424 669374
rect -23188 669138 607112 669374
rect 607348 669138 607432 669374
rect 607668 669138 607700 669374
rect -23776 669106 607700 669138
rect -23776 665974 607700 666006
rect -23776 665738 -20634 665974
rect -20398 665738 -20314 665974
rect -20078 665738 604002 665974
rect 604238 665738 604322 665974
rect 604558 665738 607700 665974
rect -23776 665654 607700 665738
rect -23776 665418 -20634 665654
rect -20398 665418 -20314 665654
rect -20078 665418 604002 665654
rect 604238 665418 604322 665654
rect 604558 665418 607700 665654
rect -23776 665386 607700 665418
rect -23776 662254 607700 662286
rect -23776 662018 -17524 662254
rect -17288 662018 -17204 662254
rect -16968 662018 580626 662254
rect 580862 662018 580946 662254
rect 581182 662018 600892 662254
rect 601128 662018 601212 662254
rect 601448 662018 607700 662254
rect -23776 661934 607700 662018
rect -23776 661698 -17524 661934
rect -17288 661698 -17204 661934
rect -16968 661698 580626 661934
rect 580862 661698 580946 661934
rect 581182 661698 600892 661934
rect 601128 661698 601212 661934
rect 601448 661698 607700 661934
rect -23776 661666 607700 661698
rect -23776 658534 607700 658566
rect -23776 658298 -14414 658534
rect -14178 658298 -14094 658534
rect -13858 658298 597782 658534
rect 598018 658298 598102 658534
rect 598338 658298 607700 658534
rect -23776 658214 607700 658298
rect -23776 657978 -14414 658214
rect -14178 657978 -14094 658214
rect -13858 657978 597782 658214
rect 598018 657978 598102 658214
rect 598338 657978 607700 658214
rect -23776 657946 607700 657978
rect -23776 654814 607700 654846
rect -23776 654578 -11304 654814
rect -11068 654578 -10984 654814
rect -10748 654578 594672 654814
rect 594908 654578 594992 654814
rect 595228 654578 607700 654814
rect -23776 654494 607700 654578
rect -23776 654258 -11304 654494
rect -11068 654258 -10984 654494
rect -10748 654258 594672 654494
rect 594908 654258 594992 654494
rect 595228 654258 607700 654494
rect -23776 654226 607700 654258
rect -23776 651094 607700 651126
rect -23776 650858 -8194 651094
rect -7958 650858 -7874 651094
rect -7638 650858 591562 651094
rect 591798 650858 591882 651094
rect 592118 650858 607700 651094
rect -23776 650774 607700 650858
rect -23776 650538 -8194 650774
rect -7958 650538 -7874 650774
rect -7638 650538 591562 650774
rect 591798 650538 591882 650774
rect 592118 650538 607700 650774
rect -23776 650506 607700 650538
rect -23776 647374 607700 647406
rect -23776 647138 -5084 647374
rect -4848 647138 -4764 647374
rect -4528 647138 7876 647374
rect 8112 647138 8196 647374
rect 8432 647138 38032 647374
rect 38268 647138 38352 647374
rect 38588 647138 74032 647374
rect 74268 647138 74352 647374
rect 74588 647138 110032 647374
rect 110268 647138 110352 647374
rect 110588 647138 146032 647374
rect 146268 647138 146352 647374
rect 146588 647138 182032 647374
rect 182268 647138 182352 647374
rect 182588 647138 218032 647374
rect 218268 647138 218352 647374
rect 218588 647138 254032 647374
rect 254268 647138 254352 647374
rect 254588 647138 290032 647374
rect 290268 647138 290352 647374
rect 290588 647138 326032 647374
rect 326268 647138 326352 647374
rect 326588 647138 362032 647374
rect 362268 647138 362352 647374
rect 362588 647138 398032 647374
rect 398268 647138 398352 647374
rect 398588 647138 434032 647374
rect 434268 647138 434352 647374
rect 434588 647138 470032 647374
rect 470268 647138 470352 647374
rect 470588 647138 506032 647374
rect 506268 647138 506352 647374
rect 506588 647138 542032 647374
rect 542268 647138 542352 647374
rect 542588 647138 571532 647374
rect 571768 647138 571852 647374
rect 572088 647138 588452 647374
rect 588688 647138 588772 647374
rect 589008 647138 607700 647374
rect -23776 647054 607700 647138
rect -23776 646818 -5084 647054
rect -4848 646818 -4764 647054
rect -4528 646818 7876 647054
rect 8112 646818 8196 647054
rect 8432 646818 38032 647054
rect 38268 646818 38352 647054
rect 38588 646818 74032 647054
rect 74268 646818 74352 647054
rect 74588 646818 110032 647054
rect 110268 646818 110352 647054
rect 110588 646818 146032 647054
rect 146268 646818 146352 647054
rect 146588 646818 182032 647054
rect 182268 646818 182352 647054
rect 182588 646818 218032 647054
rect 218268 646818 218352 647054
rect 218588 646818 254032 647054
rect 254268 646818 254352 647054
rect 254588 646818 290032 647054
rect 290268 646818 290352 647054
rect 290588 646818 326032 647054
rect 326268 646818 326352 647054
rect 326588 646818 362032 647054
rect 362268 646818 362352 647054
rect 362588 646818 398032 647054
rect 398268 646818 398352 647054
rect 398588 646818 434032 647054
rect 434268 646818 434352 647054
rect 434588 646818 470032 647054
rect 470268 646818 470352 647054
rect 470588 646818 506032 647054
rect 506268 646818 506352 647054
rect 506588 646818 542032 647054
rect 542268 646818 542352 647054
rect 542588 646818 571532 647054
rect 571768 646818 571852 647054
rect 572088 646818 588452 647054
rect 588688 646818 588772 647054
rect 589008 646818 607700 647054
rect -23776 646786 607700 646818
rect -23776 643654 607700 643686
rect -23776 643418 -1974 643654
rect -1738 643418 -1654 643654
rect -1418 643418 9116 643654
rect 9352 643418 9436 643654
rect 9672 643418 56652 643654
rect 56888 643418 56972 643654
rect 57208 643418 92652 643654
rect 92888 643418 92972 643654
rect 93208 643418 128652 643654
rect 128888 643418 128972 643654
rect 129208 643418 164652 643654
rect 164888 643418 164972 643654
rect 165208 643418 200652 643654
rect 200888 643418 200972 643654
rect 201208 643418 236652 643654
rect 236888 643418 236972 643654
rect 237208 643418 272652 643654
rect 272888 643418 272972 643654
rect 273208 643418 308652 643654
rect 308888 643418 308972 643654
rect 309208 643418 344652 643654
rect 344888 643418 344972 643654
rect 345208 643418 380652 643654
rect 380888 643418 380972 643654
rect 381208 643418 416652 643654
rect 416888 643418 416972 643654
rect 417208 643418 452652 643654
rect 452888 643418 452972 643654
rect 453208 643418 488652 643654
rect 488888 643418 488972 643654
rect 489208 643418 524652 643654
rect 524888 643418 524972 643654
rect 525208 643418 560652 643654
rect 560888 643418 560972 643654
rect 561208 643418 570292 643654
rect 570528 643418 570612 643654
rect 570848 643418 585342 643654
rect 585578 643418 585662 643654
rect 585898 643418 607700 643654
rect -23776 643334 607700 643418
rect -23776 643098 -1974 643334
rect -1738 643098 -1654 643334
rect -1418 643098 9116 643334
rect 9352 643098 9436 643334
rect 9672 643098 56652 643334
rect 56888 643098 56972 643334
rect 57208 643098 92652 643334
rect 92888 643098 92972 643334
rect 93208 643098 128652 643334
rect 128888 643098 128972 643334
rect 129208 643098 164652 643334
rect 164888 643098 164972 643334
rect 165208 643098 200652 643334
rect 200888 643098 200972 643334
rect 201208 643098 236652 643334
rect 236888 643098 236972 643334
rect 237208 643098 272652 643334
rect 272888 643098 272972 643334
rect 273208 643098 308652 643334
rect 308888 643098 308972 643334
rect 309208 643098 344652 643334
rect 344888 643098 344972 643334
rect 345208 643098 380652 643334
rect 380888 643098 380972 643334
rect 381208 643098 416652 643334
rect 416888 643098 416972 643334
rect 417208 643098 452652 643334
rect 452888 643098 452972 643334
rect 453208 643098 488652 643334
rect 488888 643098 488972 643334
rect 489208 643098 524652 643334
rect 524888 643098 524972 643334
rect 525208 643098 560652 643334
rect 560888 643098 560972 643334
rect 561208 643098 570292 643334
rect 570528 643098 570612 643334
rect 570848 643098 585342 643334
rect 585578 643098 585662 643334
rect 585898 643098 607700 643334
rect -23776 643066 607700 643098
rect -23776 629694 607700 629726
rect -23776 629458 -23744 629694
rect -23508 629458 -23424 629694
rect -23188 629458 607112 629694
rect 607348 629458 607432 629694
rect 607668 629458 607700 629694
rect -23776 629374 607700 629458
rect -23776 629138 -23744 629374
rect -23508 629138 -23424 629374
rect -23188 629138 607112 629374
rect 607348 629138 607432 629374
rect 607668 629138 607700 629374
rect -23776 629106 607700 629138
rect -23776 625974 607700 626006
rect -23776 625738 -20634 625974
rect -20398 625738 -20314 625974
rect -20078 625738 604002 625974
rect 604238 625738 604322 625974
rect 604558 625738 607700 625974
rect -23776 625654 607700 625738
rect -23776 625418 -20634 625654
rect -20398 625418 -20314 625654
rect -20078 625418 604002 625654
rect 604238 625418 604322 625654
rect 604558 625418 607700 625654
rect -23776 625386 607700 625418
rect -23776 622254 607700 622286
rect -23776 622018 -17524 622254
rect -17288 622018 -17204 622254
rect -16968 622018 580626 622254
rect 580862 622018 580946 622254
rect 581182 622018 600892 622254
rect 601128 622018 601212 622254
rect 601448 622018 607700 622254
rect -23776 621934 607700 622018
rect -23776 621698 -17524 621934
rect -17288 621698 -17204 621934
rect -16968 621698 580626 621934
rect 580862 621698 580946 621934
rect 581182 621698 600892 621934
rect 601128 621698 601212 621934
rect 601448 621698 607700 621934
rect -23776 621666 607700 621698
rect -23776 618534 607700 618566
rect -23776 618298 -14414 618534
rect -14178 618298 -14094 618534
rect -13858 618298 597782 618534
rect 598018 618298 598102 618534
rect 598338 618298 607700 618534
rect -23776 618214 607700 618298
rect -23776 617978 -14414 618214
rect -14178 617978 -14094 618214
rect -13858 617978 597782 618214
rect 598018 617978 598102 618214
rect 598338 617978 607700 618214
rect -23776 617946 607700 617978
rect -23776 614814 607700 614846
rect -23776 614578 -11304 614814
rect -11068 614578 -10984 614814
rect -10748 614578 594672 614814
rect 594908 614578 594992 614814
rect 595228 614578 607700 614814
rect -23776 614494 607700 614578
rect -23776 614258 -11304 614494
rect -11068 614258 -10984 614494
rect -10748 614258 594672 614494
rect 594908 614258 594992 614494
rect 595228 614258 607700 614494
rect -23776 614226 607700 614258
rect -23776 611094 607700 611126
rect -23776 610858 -8194 611094
rect -7958 610858 -7874 611094
rect -7638 610858 591562 611094
rect 591798 610858 591882 611094
rect 592118 610858 607700 611094
rect -23776 610774 607700 610858
rect -23776 610538 -8194 610774
rect -7958 610538 -7874 610774
rect -7638 610538 591562 610774
rect 591798 610538 591882 610774
rect 592118 610538 607700 610774
rect -23776 610506 607700 610538
rect -23776 607374 607700 607406
rect -23776 607138 -5084 607374
rect -4848 607138 -4764 607374
rect -4528 607138 7876 607374
rect 8112 607138 8196 607374
rect 8432 607138 38032 607374
rect 38268 607138 38352 607374
rect 38588 607138 74032 607374
rect 74268 607138 74352 607374
rect 74588 607138 110032 607374
rect 110268 607138 110352 607374
rect 110588 607138 146032 607374
rect 146268 607138 146352 607374
rect 146588 607138 182032 607374
rect 182268 607138 182352 607374
rect 182588 607138 218032 607374
rect 218268 607138 218352 607374
rect 218588 607138 254032 607374
rect 254268 607138 254352 607374
rect 254588 607138 290032 607374
rect 290268 607138 290352 607374
rect 290588 607138 326032 607374
rect 326268 607138 326352 607374
rect 326588 607138 362032 607374
rect 362268 607138 362352 607374
rect 362588 607138 398032 607374
rect 398268 607138 398352 607374
rect 398588 607138 434032 607374
rect 434268 607138 434352 607374
rect 434588 607138 470032 607374
rect 470268 607138 470352 607374
rect 470588 607138 506032 607374
rect 506268 607138 506352 607374
rect 506588 607138 542032 607374
rect 542268 607138 542352 607374
rect 542588 607138 571532 607374
rect 571768 607138 571852 607374
rect 572088 607138 588452 607374
rect 588688 607138 588772 607374
rect 589008 607138 607700 607374
rect -23776 607054 607700 607138
rect -23776 606818 -5084 607054
rect -4848 606818 -4764 607054
rect -4528 606818 7876 607054
rect 8112 606818 8196 607054
rect 8432 606818 38032 607054
rect 38268 606818 38352 607054
rect 38588 606818 74032 607054
rect 74268 606818 74352 607054
rect 74588 606818 110032 607054
rect 110268 606818 110352 607054
rect 110588 606818 146032 607054
rect 146268 606818 146352 607054
rect 146588 606818 182032 607054
rect 182268 606818 182352 607054
rect 182588 606818 218032 607054
rect 218268 606818 218352 607054
rect 218588 606818 254032 607054
rect 254268 606818 254352 607054
rect 254588 606818 290032 607054
rect 290268 606818 290352 607054
rect 290588 606818 326032 607054
rect 326268 606818 326352 607054
rect 326588 606818 362032 607054
rect 362268 606818 362352 607054
rect 362588 606818 398032 607054
rect 398268 606818 398352 607054
rect 398588 606818 434032 607054
rect 434268 606818 434352 607054
rect 434588 606818 470032 607054
rect 470268 606818 470352 607054
rect 470588 606818 506032 607054
rect 506268 606818 506352 607054
rect 506588 606818 542032 607054
rect 542268 606818 542352 607054
rect 542588 606818 571532 607054
rect 571768 606818 571852 607054
rect 572088 606818 588452 607054
rect 588688 606818 588772 607054
rect 589008 606818 607700 607054
rect -23776 606786 607700 606818
rect -23776 603654 607700 603686
rect -23776 603418 -1974 603654
rect -1738 603418 -1654 603654
rect -1418 603418 9116 603654
rect 9352 603418 9436 603654
rect 9672 603418 56652 603654
rect 56888 603418 56972 603654
rect 57208 603418 92652 603654
rect 92888 603418 92972 603654
rect 93208 603418 128652 603654
rect 128888 603418 128972 603654
rect 129208 603418 164652 603654
rect 164888 603418 164972 603654
rect 165208 603418 200652 603654
rect 200888 603418 200972 603654
rect 201208 603418 236652 603654
rect 236888 603418 236972 603654
rect 237208 603418 272652 603654
rect 272888 603418 272972 603654
rect 273208 603418 308652 603654
rect 308888 603418 308972 603654
rect 309208 603418 344652 603654
rect 344888 603418 344972 603654
rect 345208 603418 380652 603654
rect 380888 603418 380972 603654
rect 381208 603418 416652 603654
rect 416888 603418 416972 603654
rect 417208 603418 452652 603654
rect 452888 603418 452972 603654
rect 453208 603418 488652 603654
rect 488888 603418 488972 603654
rect 489208 603418 524652 603654
rect 524888 603418 524972 603654
rect 525208 603418 560652 603654
rect 560888 603418 560972 603654
rect 561208 603418 570292 603654
rect 570528 603418 570612 603654
rect 570848 603418 585342 603654
rect 585578 603418 585662 603654
rect 585898 603418 607700 603654
rect -23776 603334 607700 603418
rect -23776 603098 -1974 603334
rect -1738 603098 -1654 603334
rect -1418 603098 9116 603334
rect 9352 603098 9436 603334
rect 9672 603098 56652 603334
rect 56888 603098 56972 603334
rect 57208 603098 92652 603334
rect 92888 603098 92972 603334
rect 93208 603098 128652 603334
rect 128888 603098 128972 603334
rect 129208 603098 164652 603334
rect 164888 603098 164972 603334
rect 165208 603098 200652 603334
rect 200888 603098 200972 603334
rect 201208 603098 236652 603334
rect 236888 603098 236972 603334
rect 237208 603098 272652 603334
rect 272888 603098 272972 603334
rect 273208 603098 308652 603334
rect 308888 603098 308972 603334
rect 309208 603098 344652 603334
rect 344888 603098 344972 603334
rect 345208 603098 380652 603334
rect 380888 603098 380972 603334
rect 381208 603098 416652 603334
rect 416888 603098 416972 603334
rect 417208 603098 452652 603334
rect 452888 603098 452972 603334
rect 453208 603098 488652 603334
rect 488888 603098 488972 603334
rect 489208 603098 524652 603334
rect 524888 603098 524972 603334
rect 525208 603098 560652 603334
rect 560888 603098 560972 603334
rect 561208 603098 570292 603334
rect 570528 603098 570612 603334
rect 570848 603098 585342 603334
rect 585578 603098 585662 603334
rect 585898 603098 607700 603334
rect -23776 603066 607700 603098
rect -23776 589694 607700 589726
rect -23776 589458 -23744 589694
rect -23508 589458 -23424 589694
rect -23188 589458 607112 589694
rect 607348 589458 607432 589694
rect 607668 589458 607700 589694
rect -23776 589374 607700 589458
rect -23776 589138 -23744 589374
rect -23508 589138 -23424 589374
rect -23188 589138 607112 589374
rect 607348 589138 607432 589374
rect 607668 589138 607700 589374
rect -23776 589106 607700 589138
rect -23776 585974 607700 586006
rect -23776 585738 -20634 585974
rect -20398 585738 -20314 585974
rect -20078 585738 604002 585974
rect 604238 585738 604322 585974
rect 604558 585738 607700 585974
rect -23776 585654 607700 585738
rect -23776 585418 -20634 585654
rect -20398 585418 -20314 585654
rect -20078 585418 604002 585654
rect 604238 585418 604322 585654
rect 604558 585418 607700 585654
rect -23776 585386 607700 585418
rect -23776 582254 607700 582286
rect -23776 582018 -17524 582254
rect -17288 582018 -17204 582254
rect -16968 582018 580626 582254
rect 580862 582018 580946 582254
rect 581182 582018 600892 582254
rect 601128 582018 601212 582254
rect 601448 582018 607700 582254
rect -23776 581934 607700 582018
rect -23776 581698 -17524 581934
rect -17288 581698 -17204 581934
rect -16968 581698 580626 581934
rect 580862 581698 580946 581934
rect 581182 581698 600892 581934
rect 601128 581698 601212 581934
rect 601448 581698 607700 581934
rect -23776 581666 607700 581698
rect -23776 578534 607700 578566
rect -23776 578298 -14414 578534
rect -14178 578298 -14094 578534
rect -13858 578298 597782 578534
rect 598018 578298 598102 578534
rect 598338 578298 607700 578534
rect -23776 578214 607700 578298
rect -23776 577978 -14414 578214
rect -14178 577978 -14094 578214
rect -13858 577978 597782 578214
rect 598018 577978 598102 578214
rect 598338 577978 607700 578214
rect -23776 577946 607700 577978
rect -23776 574814 607700 574846
rect -23776 574578 -11304 574814
rect -11068 574578 -10984 574814
rect -10748 574578 594672 574814
rect 594908 574578 594992 574814
rect 595228 574578 607700 574814
rect -23776 574494 607700 574578
rect -23776 574258 -11304 574494
rect -11068 574258 -10984 574494
rect -10748 574258 594672 574494
rect 594908 574258 594992 574494
rect 595228 574258 607700 574494
rect -23776 574226 607700 574258
rect -23776 571094 607700 571126
rect -23776 570858 -8194 571094
rect -7958 570858 -7874 571094
rect -7638 570858 591562 571094
rect 591798 570858 591882 571094
rect 592118 570858 607700 571094
rect -23776 570774 607700 570858
rect -23776 570538 -8194 570774
rect -7958 570538 -7874 570774
rect -7638 570538 591562 570774
rect 591798 570538 591882 570774
rect 592118 570538 607700 570774
rect -23776 570506 607700 570538
rect -23776 567374 607700 567406
rect -23776 567138 -5084 567374
rect -4848 567138 -4764 567374
rect -4528 567138 7876 567374
rect 8112 567138 8196 567374
rect 8432 567138 38032 567374
rect 38268 567138 38352 567374
rect 38588 567138 74032 567374
rect 74268 567138 74352 567374
rect 74588 567138 110032 567374
rect 110268 567138 110352 567374
rect 110588 567138 146032 567374
rect 146268 567138 146352 567374
rect 146588 567138 182032 567374
rect 182268 567138 182352 567374
rect 182588 567138 218032 567374
rect 218268 567138 218352 567374
rect 218588 567138 254032 567374
rect 254268 567138 254352 567374
rect 254588 567138 290032 567374
rect 290268 567138 290352 567374
rect 290588 567138 326032 567374
rect 326268 567138 326352 567374
rect 326588 567138 362032 567374
rect 362268 567138 362352 567374
rect 362588 567138 398032 567374
rect 398268 567138 398352 567374
rect 398588 567138 434032 567374
rect 434268 567138 434352 567374
rect 434588 567138 470032 567374
rect 470268 567138 470352 567374
rect 470588 567138 506032 567374
rect 506268 567138 506352 567374
rect 506588 567138 542032 567374
rect 542268 567138 542352 567374
rect 542588 567138 571532 567374
rect 571768 567138 571852 567374
rect 572088 567138 588452 567374
rect 588688 567138 588772 567374
rect 589008 567138 607700 567374
rect -23776 567054 607700 567138
rect -23776 566818 -5084 567054
rect -4848 566818 -4764 567054
rect -4528 566818 7876 567054
rect 8112 566818 8196 567054
rect 8432 566818 38032 567054
rect 38268 566818 38352 567054
rect 38588 566818 74032 567054
rect 74268 566818 74352 567054
rect 74588 566818 110032 567054
rect 110268 566818 110352 567054
rect 110588 566818 146032 567054
rect 146268 566818 146352 567054
rect 146588 566818 182032 567054
rect 182268 566818 182352 567054
rect 182588 566818 218032 567054
rect 218268 566818 218352 567054
rect 218588 566818 254032 567054
rect 254268 566818 254352 567054
rect 254588 566818 290032 567054
rect 290268 566818 290352 567054
rect 290588 566818 326032 567054
rect 326268 566818 326352 567054
rect 326588 566818 362032 567054
rect 362268 566818 362352 567054
rect 362588 566818 398032 567054
rect 398268 566818 398352 567054
rect 398588 566818 434032 567054
rect 434268 566818 434352 567054
rect 434588 566818 470032 567054
rect 470268 566818 470352 567054
rect 470588 566818 506032 567054
rect 506268 566818 506352 567054
rect 506588 566818 542032 567054
rect 542268 566818 542352 567054
rect 542588 566818 571532 567054
rect 571768 566818 571852 567054
rect 572088 566818 588452 567054
rect 588688 566818 588772 567054
rect 589008 566818 607700 567054
rect -23776 566786 607700 566818
rect -23776 563654 607700 563686
rect -23776 563418 -1974 563654
rect -1738 563418 -1654 563654
rect -1418 563418 9116 563654
rect 9352 563418 9436 563654
rect 9672 563418 56652 563654
rect 56888 563418 56972 563654
rect 57208 563418 92652 563654
rect 92888 563418 92972 563654
rect 93208 563418 128652 563654
rect 128888 563418 128972 563654
rect 129208 563418 164652 563654
rect 164888 563418 164972 563654
rect 165208 563418 200652 563654
rect 200888 563418 200972 563654
rect 201208 563418 236652 563654
rect 236888 563418 236972 563654
rect 237208 563418 272652 563654
rect 272888 563418 272972 563654
rect 273208 563418 308652 563654
rect 308888 563418 308972 563654
rect 309208 563418 344652 563654
rect 344888 563418 344972 563654
rect 345208 563418 380652 563654
rect 380888 563418 380972 563654
rect 381208 563418 416652 563654
rect 416888 563418 416972 563654
rect 417208 563418 452652 563654
rect 452888 563418 452972 563654
rect 453208 563418 488652 563654
rect 488888 563418 488972 563654
rect 489208 563418 524652 563654
rect 524888 563418 524972 563654
rect 525208 563418 560652 563654
rect 560888 563418 560972 563654
rect 561208 563418 570292 563654
rect 570528 563418 570612 563654
rect 570848 563418 585342 563654
rect 585578 563418 585662 563654
rect 585898 563418 607700 563654
rect -23776 563334 607700 563418
rect -23776 563098 -1974 563334
rect -1738 563098 -1654 563334
rect -1418 563098 9116 563334
rect 9352 563098 9436 563334
rect 9672 563098 56652 563334
rect 56888 563098 56972 563334
rect 57208 563098 92652 563334
rect 92888 563098 92972 563334
rect 93208 563098 128652 563334
rect 128888 563098 128972 563334
rect 129208 563098 164652 563334
rect 164888 563098 164972 563334
rect 165208 563098 200652 563334
rect 200888 563098 200972 563334
rect 201208 563098 236652 563334
rect 236888 563098 236972 563334
rect 237208 563098 272652 563334
rect 272888 563098 272972 563334
rect 273208 563098 308652 563334
rect 308888 563098 308972 563334
rect 309208 563098 344652 563334
rect 344888 563098 344972 563334
rect 345208 563098 380652 563334
rect 380888 563098 380972 563334
rect 381208 563098 416652 563334
rect 416888 563098 416972 563334
rect 417208 563098 452652 563334
rect 452888 563098 452972 563334
rect 453208 563098 488652 563334
rect 488888 563098 488972 563334
rect 489208 563098 524652 563334
rect 524888 563098 524972 563334
rect 525208 563098 560652 563334
rect 560888 563098 560972 563334
rect 561208 563098 570292 563334
rect 570528 563098 570612 563334
rect 570848 563098 585342 563334
rect 585578 563098 585662 563334
rect 585898 563098 607700 563334
rect -23776 563066 607700 563098
rect -23776 549694 607700 549726
rect -23776 549458 -23744 549694
rect -23508 549458 -23424 549694
rect -23188 549458 607112 549694
rect 607348 549458 607432 549694
rect 607668 549458 607700 549694
rect -23776 549374 607700 549458
rect -23776 549138 -23744 549374
rect -23508 549138 -23424 549374
rect -23188 549138 607112 549374
rect 607348 549138 607432 549374
rect 607668 549138 607700 549374
rect -23776 549106 607700 549138
rect -23776 545974 607700 546006
rect -23776 545738 -20634 545974
rect -20398 545738 -20314 545974
rect -20078 545738 604002 545974
rect 604238 545738 604322 545974
rect 604558 545738 607700 545974
rect -23776 545654 607700 545738
rect -23776 545418 -20634 545654
rect -20398 545418 -20314 545654
rect -20078 545418 604002 545654
rect 604238 545418 604322 545654
rect 604558 545418 607700 545654
rect -23776 545386 607700 545418
rect -23776 542254 607700 542286
rect -23776 542018 -17524 542254
rect -17288 542018 -17204 542254
rect -16968 542018 580626 542254
rect 580862 542018 580946 542254
rect 581182 542018 600892 542254
rect 601128 542018 601212 542254
rect 601448 542018 607700 542254
rect -23776 541934 607700 542018
rect -23776 541698 -17524 541934
rect -17288 541698 -17204 541934
rect -16968 541698 580626 541934
rect 580862 541698 580946 541934
rect 581182 541698 600892 541934
rect 601128 541698 601212 541934
rect 601448 541698 607700 541934
rect -23776 541666 607700 541698
rect -23776 538534 607700 538566
rect -23776 538298 -14414 538534
rect -14178 538298 -14094 538534
rect -13858 538298 597782 538534
rect 598018 538298 598102 538534
rect 598338 538298 607700 538534
rect -23776 538214 607700 538298
rect -23776 537978 -14414 538214
rect -14178 537978 -14094 538214
rect -13858 537978 597782 538214
rect 598018 537978 598102 538214
rect 598338 537978 607700 538214
rect -23776 537946 607700 537978
rect -23776 534814 607700 534846
rect -23776 534578 -11304 534814
rect -11068 534578 -10984 534814
rect -10748 534578 594672 534814
rect 594908 534578 594992 534814
rect 595228 534578 607700 534814
rect -23776 534494 607700 534578
rect -23776 534258 -11304 534494
rect -11068 534258 -10984 534494
rect -10748 534258 594672 534494
rect 594908 534258 594992 534494
rect 595228 534258 607700 534494
rect -23776 534226 607700 534258
rect -23776 531094 607700 531126
rect -23776 530858 -8194 531094
rect -7958 530858 -7874 531094
rect -7638 530858 591562 531094
rect 591798 530858 591882 531094
rect 592118 530858 607700 531094
rect -23776 530774 607700 530858
rect -23776 530538 -8194 530774
rect -7958 530538 -7874 530774
rect -7638 530538 591562 530774
rect 591798 530538 591882 530774
rect 592118 530538 607700 530774
rect -23776 530506 607700 530538
rect -23776 527374 607700 527406
rect -23776 527138 -5084 527374
rect -4848 527138 -4764 527374
rect -4528 527138 7876 527374
rect 8112 527138 8196 527374
rect 8432 527138 38032 527374
rect 38268 527138 38352 527374
rect 38588 527138 74032 527374
rect 74268 527138 74352 527374
rect 74588 527138 110032 527374
rect 110268 527138 110352 527374
rect 110588 527138 146032 527374
rect 146268 527138 146352 527374
rect 146588 527138 182032 527374
rect 182268 527138 182352 527374
rect 182588 527138 218032 527374
rect 218268 527138 218352 527374
rect 218588 527138 254032 527374
rect 254268 527138 254352 527374
rect 254588 527138 290032 527374
rect 290268 527138 290352 527374
rect 290588 527138 326032 527374
rect 326268 527138 326352 527374
rect 326588 527138 362032 527374
rect 362268 527138 362352 527374
rect 362588 527138 398032 527374
rect 398268 527138 398352 527374
rect 398588 527138 434032 527374
rect 434268 527138 434352 527374
rect 434588 527138 470032 527374
rect 470268 527138 470352 527374
rect 470588 527138 506032 527374
rect 506268 527138 506352 527374
rect 506588 527138 542032 527374
rect 542268 527138 542352 527374
rect 542588 527138 571532 527374
rect 571768 527138 571852 527374
rect 572088 527138 588452 527374
rect 588688 527138 588772 527374
rect 589008 527138 607700 527374
rect -23776 527054 607700 527138
rect -23776 526818 -5084 527054
rect -4848 526818 -4764 527054
rect -4528 526818 7876 527054
rect 8112 526818 8196 527054
rect 8432 526818 38032 527054
rect 38268 526818 38352 527054
rect 38588 526818 74032 527054
rect 74268 526818 74352 527054
rect 74588 526818 110032 527054
rect 110268 526818 110352 527054
rect 110588 526818 146032 527054
rect 146268 526818 146352 527054
rect 146588 526818 182032 527054
rect 182268 526818 182352 527054
rect 182588 526818 218032 527054
rect 218268 526818 218352 527054
rect 218588 526818 254032 527054
rect 254268 526818 254352 527054
rect 254588 526818 290032 527054
rect 290268 526818 290352 527054
rect 290588 526818 326032 527054
rect 326268 526818 326352 527054
rect 326588 526818 362032 527054
rect 362268 526818 362352 527054
rect 362588 526818 398032 527054
rect 398268 526818 398352 527054
rect 398588 526818 434032 527054
rect 434268 526818 434352 527054
rect 434588 526818 470032 527054
rect 470268 526818 470352 527054
rect 470588 526818 506032 527054
rect 506268 526818 506352 527054
rect 506588 526818 542032 527054
rect 542268 526818 542352 527054
rect 542588 526818 571532 527054
rect 571768 526818 571852 527054
rect 572088 526818 588452 527054
rect 588688 526818 588772 527054
rect 589008 526818 607700 527054
rect -23776 526786 607700 526818
rect -23776 523654 607700 523686
rect -23776 523418 -1974 523654
rect -1738 523418 -1654 523654
rect -1418 523418 9116 523654
rect 9352 523418 9436 523654
rect 9672 523418 56652 523654
rect 56888 523418 56972 523654
rect 57208 523418 92652 523654
rect 92888 523418 92972 523654
rect 93208 523418 128652 523654
rect 128888 523418 128972 523654
rect 129208 523418 164652 523654
rect 164888 523418 164972 523654
rect 165208 523418 200652 523654
rect 200888 523418 200972 523654
rect 201208 523418 236652 523654
rect 236888 523418 236972 523654
rect 237208 523418 272652 523654
rect 272888 523418 272972 523654
rect 273208 523418 308652 523654
rect 308888 523418 308972 523654
rect 309208 523418 344652 523654
rect 344888 523418 344972 523654
rect 345208 523418 380652 523654
rect 380888 523418 380972 523654
rect 381208 523418 416652 523654
rect 416888 523418 416972 523654
rect 417208 523418 452652 523654
rect 452888 523418 452972 523654
rect 453208 523418 488652 523654
rect 488888 523418 488972 523654
rect 489208 523418 524652 523654
rect 524888 523418 524972 523654
rect 525208 523418 560652 523654
rect 560888 523418 560972 523654
rect 561208 523418 570292 523654
rect 570528 523418 570612 523654
rect 570848 523418 585342 523654
rect 585578 523418 585662 523654
rect 585898 523418 607700 523654
rect -23776 523334 607700 523418
rect -23776 523098 -1974 523334
rect -1738 523098 -1654 523334
rect -1418 523098 9116 523334
rect 9352 523098 9436 523334
rect 9672 523098 56652 523334
rect 56888 523098 56972 523334
rect 57208 523098 92652 523334
rect 92888 523098 92972 523334
rect 93208 523098 128652 523334
rect 128888 523098 128972 523334
rect 129208 523098 164652 523334
rect 164888 523098 164972 523334
rect 165208 523098 200652 523334
rect 200888 523098 200972 523334
rect 201208 523098 236652 523334
rect 236888 523098 236972 523334
rect 237208 523098 272652 523334
rect 272888 523098 272972 523334
rect 273208 523098 308652 523334
rect 308888 523098 308972 523334
rect 309208 523098 344652 523334
rect 344888 523098 344972 523334
rect 345208 523098 380652 523334
rect 380888 523098 380972 523334
rect 381208 523098 416652 523334
rect 416888 523098 416972 523334
rect 417208 523098 452652 523334
rect 452888 523098 452972 523334
rect 453208 523098 488652 523334
rect 488888 523098 488972 523334
rect 489208 523098 524652 523334
rect 524888 523098 524972 523334
rect 525208 523098 560652 523334
rect 560888 523098 560972 523334
rect 561208 523098 570292 523334
rect 570528 523098 570612 523334
rect 570848 523098 585342 523334
rect 585578 523098 585662 523334
rect 585898 523098 607700 523334
rect -23776 523066 607700 523098
rect -23776 509694 607700 509726
rect -23776 509458 -23744 509694
rect -23508 509458 -23424 509694
rect -23188 509458 607112 509694
rect 607348 509458 607432 509694
rect 607668 509458 607700 509694
rect -23776 509374 607700 509458
rect -23776 509138 -23744 509374
rect -23508 509138 -23424 509374
rect -23188 509138 607112 509374
rect 607348 509138 607432 509374
rect 607668 509138 607700 509374
rect -23776 509106 607700 509138
rect -23776 505974 607700 506006
rect -23776 505738 -20634 505974
rect -20398 505738 -20314 505974
rect -20078 505738 604002 505974
rect 604238 505738 604322 505974
rect 604558 505738 607700 505974
rect -23776 505654 607700 505738
rect -23776 505418 -20634 505654
rect -20398 505418 -20314 505654
rect -20078 505418 604002 505654
rect 604238 505418 604322 505654
rect 604558 505418 607700 505654
rect -23776 505386 607700 505418
rect -23776 502254 607700 502286
rect -23776 502018 -17524 502254
rect -17288 502018 -17204 502254
rect -16968 502018 580626 502254
rect 580862 502018 580946 502254
rect 581182 502018 600892 502254
rect 601128 502018 601212 502254
rect 601448 502018 607700 502254
rect -23776 501934 607700 502018
rect -23776 501698 -17524 501934
rect -17288 501698 -17204 501934
rect -16968 501698 580626 501934
rect 580862 501698 580946 501934
rect 581182 501698 600892 501934
rect 601128 501698 601212 501934
rect 601448 501698 607700 501934
rect -23776 501666 607700 501698
rect -23776 498534 607700 498566
rect -23776 498298 -14414 498534
rect -14178 498298 -14094 498534
rect -13858 498298 597782 498534
rect 598018 498298 598102 498534
rect 598338 498298 607700 498534
rect -23776 498214 607700 498298
rect -23776 497978 -14414 498214
rect -14178 497978 -14094 498214
rect -13858 497978 597782 498214
rect 598018 497978 598102 498214
rect 598338 497978 607700 498214
rect -23776 497946 607700 497978
rect -23776 494814 607700 494846
rect -23776 494578 -11304 494814
rect -11068 494578 -10984 494814
rect -10748 494578 594672 494814
rect 594908 494578 594992 494814
rect 595228 494578 607700 494814
rect -23776 494494 607700 494578
rect -23776 494258 -11304 494494
rect -11068 494258 -10984 494494
rect -10748 494258 594672 494494
rect 594908 494258 594992 494494
rect 595228 494258 607700 494494
rect -23776 494226 607700 494258
rect -23776 491094 607700 491126
rect -23776 490858 -8194 491094
rect -7958 490858 -7874 491094
rect -7638 490858 591562 491094
rect 591798 490858 591882 491094
rect 592118 490858 607700 491094
rect -23776 490774 607700 490858
rect -23776 490538 -8194 490774
rect -7958 490538 -7874 490774
rect -7638 490538 591562 490774
rect 591798 490538 591882 490774
rect 592118 490538 607700 490774
rect -23776 490506 607700 490538
rect -23776 487374 607700 487406
rect -23776 487138 -5084 487374
rect -4848 487138 -4764 487374
rect -4528 487138 7876 487374
rect 8112 487138 8196 487374
rect 8432 487138 38032 487374
rect 38268 487138 38352 487374
rect 38588 487138 60622 487374
rect 60858 487138 159098 487374
rect 159334 487138 182032 487374
rect 182268 487138 182352 487374
rect 182588 487138 185622 487374
rect 185858 487138 284098 487374
rect 284334 487138 290032 487374
rect 290268 487138 290352 487374
rect 290588 487138 310622 487374
rect 310858 487138 409098 487374
rect 409334 487138 434032 487374
rect 434268 487138 434352 487374
rect 434588 487138 436622 487374
rect 436858 487138 535098 487374
rect 535334 487138 542032 487374
rect 542268 487138 542352 487374
rect 542588 487138 571532 487374
rect 571768 487138 571852 487374
rect 572088 487138 588452 487374
rect 588688 487138 588772 487374
rect 589008 487138 607700 487374
rect -23776 487054 607700 487138
rect -23776 486818 -5084 487054
rect -4848 486818 -4764 487054
rect -4528 486818 7876 487054
rect 8112 486818 8196 487054
rect 8432 486818 38032 487054
rect 38268 486818 38352 487054
rect 38588 486818 60622 487054
rect 60858 486818 159098 487054
rect 159334 486818 182032 487054
rect 182268 486818 182352 487054
rect 182588 486818 185622 487054
rect 185858 486818 284098 487054
rect 284334 486818 290032 487054
rect 290268 486818 290352 487054
rect 290588 486818 310622 487054
rect 310858 486818 409098 487054
rect 409334 486818 434032 487054
rect 434268 486818 434352 487054
rect 434588 486818 436622 487054
rect 436858 486818 535098 487054
rect 535334 486818 542032 487054
rect 542268 486818 542352 487054
rect 542588 486818 571532 487054
rect 571768 486818 571852 487054
rect 572088 486818 588452 487054
rect 588688 486818 588772 487054
rect 589008 486818 607700 487054
rect -23776 486786 607700 486818
rect -23776 483654 607700 483686
rect -23776 483418 -1974 483654
rect -1738 483418 -1654 483654
rect -1418 483418 9116 483654
rect 9352 483418 9436 483654
rect 9672 483418 56652 483654
rect 56888 483418 56972 483654
rect 57208 483418 61342 483654
rect 61578 483418 158378 483654
rect 158614 483418 164652 483654
rect 164888 483418 164972 483654
rect 165208 483418 186342 483654
rect 186578 483418 283378 483654
rect 283614 483418 308652 483654
rect 308888 483418 308972 483654
rect 309208 483418 311342 483654
rect 311578 483418 408378 483654
rect 408614 483418 416652 483654
rect 416888 483418 416972 483654
rect 417208 483418 437342 483654
rect 437578 483418 534378 483654
rect 534614 483418 560652 483654
rect 560888 483418 560972 483654
rect 561208 483418 570292 483654
rect 570528 483418 570612 483654
rect 570848 483418 585342 483654
rect 585578 483418 585662 483654
rect 585898 483418 607700 483654
rect -23776 483334 607700 483418
rect -23776 483098 -1974 483334
rect -1738 483098 -1654 483334
rect -1418 483098 9116 483334
rect 9352 483098 9436 483334
rect 9672 483098 56652 483334
rect 56888 483098 56972 483334
rect 57208 483098 61342 483334
rect 61578 483098 158378 483334
rect 158614 483098 164652 483334
rect 164888 483098 164972 483334
rect 165208 483098 186342 483334
rect 186578 483098 283378 483334
rect 283614 483098 308652 483334
rect 308888 483098 308972 483334
rect 309208 483098 311342 483334
rect 311578 483098 408378 483334
rect 408614 483098 416652 483334
rect 416888 483098 416972 483334
rect 417208 483098 437342 483334
rect 437578 483098 534378 483334
rect 534614 483098 560652 483334
rect 560888 483098 560972 483334
rect 561208 483098 570292 483334
rect 570528 483098 570612 483334
rect 570848 483098 585342 483334
rect 585578 483098 585662 483334
rect 585898 483098 607700 483334
rect -23776 483066 607700 483098
rect -23776 469694 607700 469726
rect -23776 469458 -23744 469694
rect -23508 469458 -23424 469694
rect -23188 469458 607112 469694
rect 607348 469458 607432 469694
rect 607668 469458 607700 469694
rect -23776 469374 607700 469458
rect -23776 469138 -23744 469374
rect -23508 469138 -23424 469374
rect -23188 469138 607112 469374
rect 607348 469138 607432 469374
rect 607668 469138 607700 469374
rect -23776 469106 607700 469138
rect -23776 465974 607700 466006
rect -23776 465738 -20634 465974
rect -20398 465738 -20314 465974
rect -20078 465738 604002 465974
rect 604238 465738 604322 465974
rect 604558 465738 607700 465974
rect -23776 465654 607700 465738
rect -23776 465418 -20634 465654
rect -20398 465418 -20314 465654
rect -20078 465418 604002 465654
rect 604238 465418 604322 465654
rect 604558 465418 607700 465654
rect -23776 465386 607700 465418
rect -23776 462254 607700 462286
rect -23776 462018 -17524 462254
rect -17288 462018 -17204 462254
rect -16968 462018 580626 462254
rect 580862 462018 580946 462254
rect 581182 462018 600892 462254
rect 601128 462018 601212 462254
rect 601448 462018 607700 462254
rect -23776 461934 607700 462018
rect -23776 461698 -17524 461934
rect -17288 461698 -17204 461934
rect -16968 461698 580626 461934
rect 580862 461698 580946 461934
rect 581182 461698 600892 461934
rect 601128 461698 601212 461934
rect 601448 461698 607700 461934
rect -23776 461666 607700 461698
rect -23776 458534 607700 458566
rect -23776 458298 -14414 458534
rect -14178 458298 -14094 458534
rect -13858 458298 597782 458534
rect 598018 458298 598102 458534
rect 598338 458298 607700 458534
rect -23776 458214 607700 458298
rect -23776 457978 -14414 458214
rect -14178 457978 -14094 458214
rect -13858 457978 597782 458214
rect 598018 457978 598102 458214
rect 598338 457978 607700 458214
rect -23776 457946 607700 457978
rect -23776 454814 607700 454846
rect -23776 454578 -11304 454814
rect -11068 454578 -10984 454814
rect -10748 454578 594672 454814
rect 594908 454578 594992 454814
rect 595228 454578 607700 454814
rect -23776 454494 607700 454578
rect -23776 454258 -11304 454494
rect -11068 454258 -10984 454494
rect -10748 454258 594672 454494
rect 594908 454258 594992 454494
rect 595228 454258 607700 454494
rect -23776 454226 607700 454258
rect -23776 451094 607700 451126
rect -23776 450858 -8194 451094
rect -7958 450858 -7874 451094
rect -7638 450858 591562 451094
rect 591798 450858 591882 451094
rect 592118 450858 607700 451094
rect -23776 450774 607700 450858
rect -23776 450538 -8194 450774
rect -7958 450538 -7874 450774
rect -7638 450538 591562 450774
rect 591798 450538 591882 450774
rect 592118 450538 607700 450774
rect -23776 450506 607700 450538
rect -23776 447374 607700 447406
rect -23776 447138 -5084 447374
rect -4848 447138 -4764 447374
rect -4528 447138 7876 447374
rect 8112 447138 8196 447374
rect 8432 447138 38032 447374
rect 38268 447138 38352 447374
rect 38588 447138 60622 447374
rect 60858 447138 159098 447374
rect 159334 447138 182032 447374
rect 182268 447138 182352 447374
rect 182588 447138 185622 447374
rect 185858 447138 284098 447374
rect 284334 447138 290032 447374
rect 290268 447138 290352 447374
rect 290588 447138 310622 447374
rect 310858 447138 409098 447374
rect 409334 447138 434032 447374
rect 434268 447138 434352 447374
rect 434588 447138 436622 447374
rect 436858 447138 535098 447374
rect 535334 447138 542032 447374
rect 542268 447138 542352 447374
rect 542588 447138 571532 447374
rect 571768 447138 571852 447374
rect 572088 447138 588452 447374
rect 588688 447138 588772 447374
rect 589008 447138 607700 447374
rect -23776 447054 607700 447138
rect -23776 446818 -5084 447054
rect -4848 446818 -4764 447054
rect -4528 446818 7876 447054
rect 8112 446818 8196 447054
rect 8432 446818 38032 447054
rect 38268 446818 38352 447054
rect 38588 446818 60622 447054
rect 60858 446818 159098 447054
rect 159334 446818 182032 447054
rect 182268 446818 182352 447054
rect 182588 446818 185622 447054
rect 185858 446818 284098 447054
rect 284334 446818 290032 447054
rect 290268 446818 290352 447054
rect 290588 446818 310622 447054
rect 310858 446818 409098 447054
rect 409334 446818 434032 447054
rect 434268 446818 434352 447054
rect 434588 446818 436622 447054
rect 436858 446818 535098 447054
rect 535334 446818 542032 447054
rect 542268 446818 542352 447054
rect 542588 446818 571532 447054
rect 571768 446818 571852 447054
rect 572088 446818 588452 447054
rect 588688 446818 588772 447054
rect 589008 446818 607700 447054
rect -23776 446786 607700 446818
rect -23776 443654 607700 443686
rect -23776 443418 -1974 443654
rect -1738 443418 -1654 443654
rect -1418 443418 9116 443654
rect 9352 443418 9436 443654
rect 9672 443418 56652 443654
rect 56888 443418 56972 443654
rect 57208 443418 61342 443654
rect 61578 443418 158378 443654
rect 158614 443418 164652 443654
rect 164888 443418 164972 443654
rect 165208 443418 186342 443654
rect 186578 443418 283378 443654
rect 283614 443418 308652 443654
rect 308888 443418 308972 443654
rect 309208 443418 311342 443654
rect 311578 443418 408378 443654
rect 408614 443418 416652 443654
rect 416888 443418 416972 443654
rect 417208 443418 437342 443654
rect 437578 443418 534378 443654
rect 534614 443418 560652 443654
rect 560888 443418 560972 443654
rect 561208 443418 570292 443654
rect 570528 443418 570612 443654
rect 570848 443418 585342 443654
rect 585578 443418 585662 443654
rect 585898 443418 607700 443654
rect -23776 443334 607700 443418
rect -23776 443098 -1974 443334
rect -1738 443098 -1654 443334
rect -1418 443098 9116 443334
rect 9352 443098 9436 443334
rect 9672 443098 56652 443334
rect 56888 443098 56972 443334
rect 57208 443098 61342 443334
rect 61578 443098 158378 443334
rect 158614 443098 164652 443334
rect 164888 443098 164972 443334
rect 165208 443098 186342 443334
rect 186578 443098 283378 443334
rect 283614 443098 308652 443334
rect 308888 443098 308972 443334
rect 309208 443098 311342 443334
rect 311578 443098 408378 443334
rect 408614 443098 416652 443334
rect 416888 443098 416972 443334
rect 417208 443098 437342 443334
rect 437578 443098 534378 443334
rect 534614 443098 560652 443334
rect 560888 443098 560972 443334
rect 561208 443098 570292 443334
rect 570528 443098 570612 443334
rect 570848 443098 585342 443334
rect 585578 443098 585662 443334
rect 585898 443098 607700 443334
rect -23776 443066 607700 443098
rect 61280 433244 61640 433300
rect 61280 433008 61342 433244
rect 61578 433008 61640 433244
rect 61280 432952 61640 433008
rect 62952 433244 63300 433300
rect 62952 433008 63008 433244
rect 63244 433008 63300 433244
rect 62952 432952 63300 433008
rect 281656 433244 282004 433300
rect 281656 433008 281712 433244
rect 281948 433008 282004 433244
rect 281656 432952 282004 433008
rect 283316 433244 283676 433300
rect 283316 433008 283378 433244
rect 283614 433008 283676 433244
rect 283316 432952 283676 433008
rect 311280 433244 311640 433300
rect 311280 433008 311342 433244
rect 311578 433008 311640 433244
rect 311280 432952 311640 433008
rect 312952 433244 313300 433300
rect 312952 433008 313008 433244
rect 313244 433008 313300 433244
rect 312952 432952 313300 433008
rect 532656 433244 533004 433300
rect 532656 433008 532712 433244
rect 532948 433008 533004 433244
rect 532656 432952 533004 433008
rect 534316 433244 534676 433300
rect 534316 433008 534378 433244
rect 534614 433008 534676 433244
rect 534316 432952 534676 433008
rect 157336 432564 157684 432620
rect 157336 432328 157392 432564
rect 157628 432328 157684 432564
rect 157336 432272 157684 432328
rect 159036 432564 159396 432620
rect 159036 432328 159098 432564
rect 159334 432328 159396 432564
rect 159036 432272 159396 432328
rect 185560 432564 185920 432620
rect 185560 432328 185622 432564
rect 185858 432328 185920 432564
rect 185560 432272 185920 432328
rect 187272 432564 187620 432620
rect 187272 432328 187328 432564
rect 187564 432328 187620 432564
rect 187272 432272 187620 432328
rect 407336 432564 407684 432620
rect 407336 432328 407392 432564
rect 407628 432328 407684 432564
rect 407336 432272 407684 432328
rect 409036 432564 409396 432620
rect 409036 432328 409098 432564
rect 409334 432328 409396 432564
rect 409036 432272 409396 432328
rect 436560 432564 436920 432620
rect 436560 432328 436622 432564
rect 436858 432328 436920 432564
rect 436560 432272 436920 432328
rect 438272 432564 438620 432620
rect 438272 432328 438328 432564
rect 438564 432328 438620 432564
rect 438272 432272 438620 432328
rect -23776 429694 607700 429726
rect -23776 429458 -23744 429694
rect -23508 429458 -23424 429694
rect -23188 429458 607112 429694
rect 607348 429458 607432 429694
rect 607668 429458 607700 429694
rect -23776 429374 607700 429458
rect -23776 429138 -23744 429374
rect -23508 429138 -23424 429374
rect -23188 429138 607112 429374
rect 607348 429138 607432 429374
rect 607668 429138 607700 429374
rect -23776 429106 607700 429138
rect -23776 425974 607700 426006
rect -23776 425738 -20634 425974
rect -20398 425738 -20314 425974
rect -20078 425738 604002 425974
rect 604238 425738 604322 425974
rect 604558 425738 607700 425974
rect -23776 425654 607700 425738
rect -23776 425418 -20634 425654
rect -20398 425418 -20314 425654
rect -20078 425418 604002 425654
rect 604238 425418 604322 425654
rect 604558 425418 607700 425654
rect -23776 425386 607700 425418
rect -23776 422254 607700 422286
rect -23776 422018 -17524 422254
rect -17288 422018 -17204 422254
rect -16968 422018 580626 422254
rect 580862 422018 580946 422254
rect 581182 422018 600892 422254
rect 601128 422018 601212 422254
rect 601448 422018 607700 422254
rect -23776 421934 607700 422018
rect -23776 421698 -17524 421934
rect -17288 421698 -17204 421934
rect -16968 421698 580626 421934
rect 580862 421698 580946 421934
rect 581182 421698 600892 421934
rect 601128 421698 601212 421934
rect 601448 421698 607700 421934
rect -23776 421666 607700 421698
rect -23776 418534 607700 418566
rect -23776 418298 -14414 418534
rect -14178 418298 -14094 418534
rect -13858 418298 597782 418534
rect 598018 418298 598102 418534
rect 598338 418298 607700 418534
rect -23776 418214 607700 418298
rect -23776 417978 -14414 418214
rect -14178 417978 -14094 418214
rect -13858 417978 597782 418214
rect 598018 417978 598102 418214
rect 598338 417978 607700 418214
rect -23776 417946 607700 417978
rect -23776 414814 607700 414846
rect -23776 414578 -11304 414814
rect -11068 414578 -10984 414814
rect -10748 414578 594672 414814
rect 594908 414578 594992 414814
rect 595228 414578 607700 414814
rect -23776 414494 607700 414578
rect -23776 414258 -11304 414494
rect -11068 414258 -10984 414494
rect -10748 414258 594672 414494
rect 594908 414258 594992 414494
rect 595228 414258 607700 414494
rect -23776 414226 607700 414258
rect -23776 411094 607700 411126
rect -23776 410858 -8194 411094
rect -7958 410858 -7874 411094
rect -7638 410858 591562 411094
rect 591798 410858 591882 411094
rect 592118 410858 607700 411094
rect -23776 410774 607700 410858
rect -23776 410538 -8194 410774
rect -7958 410538 -7874 410774
rect -7638 410538 591562 410774
rect 591798 410538 591882 410774
rect 592118 410538 607700 410774
rect -23776 410506 607700 410538
rect -23776 407374 607700 407406
rect -23776 407138 -5084 407374
rect -4848 407138 -4764 407374
rect -4528 407138 7876 407374
rect 8112 407138 8196 407374
rect 8432 407138 38032 407374
rect 38268 407138 38352 407374
rect 38588 407138 74032 407374
rect 74268 407138 74352 407374
rect 74588 407138 110032 407374
rect 110268 407138 110352 407374
rect 110588 407138 146032 407374
rect 146268 407138 146352 407374
rect 146588 407138 182032 407374
rect 182268 407138 182352 407374
rect 182588 407138 218032 407374
rect 218268 407138 218352 407374
rect 218588 407138 254032 407374
rect 254268 407138 254352 407374
rect 254588 407138 290032 407374
rect 290268 407138 290352 407374
rect 290588 407138 326032 407374
rect 326268 407138 326352 407374
rect 326588 407138 362032 407374
rect 362268 407138 362352 407374
rect 362588 407138 398032 407374
rect 398268 407138 398352 407374
rect 398588 407138 434032 407374
rect 434268 407138 434352 407374
rect 434588 407138 470032 407374
rect 470268 407138 470352 407374
rect 470588 407138 506032 407374
rect 506268 407138 506352 407374
rect 506588 407138 542032 407374
rect 542268 407138 542352 407374
rect 542588 407138 571532 407374
rect 571768 407138 571852 407374
rect 572088 407138 588452 407374
rect 588688 407138 588772 407374
rect 589008 407138 607700 407374
rect -23776 407054 607700 407138
rect -23776 406818 -5084 407054
rect -4848 406818 -4764 407054
rect -4528 406818 7876 407054
rect 8112 406818 8196 407054
rect 8432 406818 38032 407054
rect 38268 406818 38352 407054
rect 38588 406818 74032 407054
rect 74268 406818 74352 407054
rect 74588 406818 110032 407054
rect 110268 406818 110352 407054
rect 110588 406818 146032 407054
rect 146268 406818 146352 407054
rect 146588 406818 182032 407054
rect 182268 406818 182352 407054
rect 182588 406818 218032 407054
rect 218268 406818 218352 407054
rect 218588 406818 254032 407054
rect 254268 406818 254352 407054
rect 254588 406818 290032 407054
rect 290268 406818 290352 407054
rect 290588 406818 326032 407054
rect 326268 406818 326352 407054
rect 326588 406818 362032 407054
rect 362268 406818 362352 407054
rect 362588 406818 398032 407054
rect 398268 406818 398352 407054
rect 398588 406818 434032 407054
rect 434268 406818 434352 407054
rect 434588 406818 470032 407054
rect 470268 406818 470352 407054
rect 470588 406818 506032 407054
rect 506268 406818 506352 407054
rect 506588 406818 542032 407054
rect 542268 406818 542352 407054
rect 542588 406818 571532 407054
rect 571768 406818 571852 407054
rect 572088 406818 588452 407054
rect 588688 406818 588772 407054
rect 589008 406818 607700 407054
rect -23776 406786 607700 406818
rect -23776 403654 607700 403686
rect -23776 403418 -1974 403654
rect -1738 403418 -1654 403654
rect -1418 403418 9116 403654
rect 9352 403418 9436 403654
rect 9672 403418 56652 403654
rect 56888 403418 56972 403654
rect 57208 403418 92652 403654
rect 92888 403418 92972 403654
rect 93208 403418 128652 403654
rect 128888 403418 128972 403654
rect 129208 403418 164652 403654
rect 164888 403418 164972 403654
rect 165208 403418 200652 403654
rect 200888 403418 200972 403654
rect 201208 403418 236652 403654
rect 236888 403418 236972 403654
rect 237208 403418 272652 403654
rect 272888 403418 272972 403654
rect 273208 403418 308652 403654
rect 308888 403418 308972 403654
rect 309208 403418 344652 403654
rect 344888 403418 344972 403654
rect 345208 403418 380652 403654
rect 380888 403418 380972 403654
rect 381208 403418 416652 403654
rect 416888 403418 416972 403654
rect 417208 403418 452652 403654
rect 452888 403418 452972 403654
rect 453208 403418 488652 403654
rect 488888 403418 488972 403654
rect 489208 403418 524652 403654
rect 524888 403418 524972 403654
rect 525208 403418 560652 403654
rect 560888 403418 560972 403654
rect 561208 403418 570292 403654
rect 570528 403418 570612 403654
rect 570848 403418 585342 403654
rect 585578 403418 585662 403654
rect 585898 403418 607700 403654
rect -23776 403334 607700 403418
rect -23776 403098 -1974 403334
rect -1738 403098 -1654 403334
rect -1418 403098 9116 403334
rect 9352 403098 9436 403334
rect 9672 403098 56652 403334
rect 56888 403098 56972 403334
rect 57208 403098 92652 403334
rect 92888 403098 92972 403334
rect 93208 403098 128652 403334
rect 128888 403098 128972 403334
rect 129208 403098 164652 403334
rect 164888 403098 164972 403334
rect 165208 403098 200652 403334
rect 200888 403098 200972 403334
rect 201208 403098 236652 403334
rect 236888 403098 236972 403334
rect 237208 403098 272652 403334
rect 272888 403098 272972 403334
rect 273208 403098 308652 403334
rect 308888 403098 308972 403334
rect 309208 403098 344652 403334
rect 344888 403098 344972 403334
rect 345208 403098 380652 403334
rect 380888 403098 380972 403334
rect 381208 403098 416652 403334
rect 416888 403098 416972 403334
rect 417208 403098 452652 403334
rect 452888 403098 452972 403334
rect 453208 403098 488652 403334
rect 488888 403098 488972 403334
rect 489208 403098 524652 403334
rect 524888 403098 524972 403334
rect 525208 403098 560652 403334
rect 560888 403098 560972 403334
rect 561208 403098 570292 403334
rect 570528 403098 570612 403334
rect 570848 403098 585342 403334
rect 585578 403098 585662 403334
rect 585898 403098 607700 403334
rect -23776 403066 607700 403098
rect -23776 389694 607700 389726
rect -23776 389458 -23744 389694
rect -23508 389458 -23424 389694
rect -23188 389458 607112 389694
rect 607348 389458 607432 389694
rect 607668 389458 607700 389694
rect -23776 389374 607700 389458
rect -23776 389138 -23744 389374
rect -23508 389138 -23424 389374
rect -23188 389138 607112 389374
rect 607348 389138 607432 389374
rect 607668 389138 607700 389374
rect -23776 389106 607700 389138
rect -23776 385974 607700 386006
rect -23776 385738 -20634 385974
rect -20398 385738 -20314 385974
rect -20078 385738 604002 385974
rect 604238 385738 604322 385974
rect 604558 385738 607700 385974
rect -23776 385654 607700 385738
rect -23776 385418 -20634 385654
rect -20398 385418 -20314 385654
rect -20078 385418 604002 385654
rect 604238 385418 604322 385654
rect 604558 385418 607700 385654
rect -23776 385386 607700 385418
rect -23776 382254 607700 382286
rect -23776 382018 -17524 382254
rect -17288 382018 -17204 382254
rect -16968 382018 580626 382254
rect 580862 382018 580946 382254
rect 581182 382018 600892 382254
rect 601128 382018 601212 382254
rect 601448 382018 607700 382254
rect -23776 381934 607700 382018
rect -23776 381698 -17524 381934
rect -17288 381698 -17204 381934
rect -16968 381698 580626 381934
rect 580862 381698 580946 381934
rect 581182 381698 600892 381934
rect 601128 381698 601212 381934
rect 601448 381698 607700 381934
rect -23776 381666 607700 381698
rect -23776 378534 607700 378566
rect -23776 378298 -14414 378534
rect -14178 378298 -14094 378534
rect -13858 378298 597782 378534
rect 598018 378298 598102 378534
rect 598338 378298 607700 378534
rect -23776 378214 607700 378298
rect -23776 377978 -14414 378214
rect -14178 377978 -14094 378214
rect -13858 377978 597782 378214
rect 598018 377978 598102 378214
rect 598338 377978 607700 378214
rect -23776 377946 607700 377978
rect -23776 374814 607700 374846
rect -23776 374578 -11304 374814
rect -11068 374578 -10984 374814
rect -10748 374578 594672 374814
rect 594908 374578 594992 374814
rect 595228 374578 607700 374814
rect -23776 374494 607700 374578
rect -23776 374258 -11304 374494
rect -11068 374258 -10984 374494
rect -10748 374258 594672 374494
rect 594908 374258 594992 374494
rect 595228 374258 607700 374494
rect -23776 374226 607700 374258
rect -23776 371094 607700 371126
rect -23776 370858 -8194 371094
rect -7958 370858 -7874 371094
rect -7638 370858 591562 371094
rect 591798 370858 591882 371094
rect 592118 370858 607700 371094
rect -23776 370774 607700 370858
rect -23776 370538 -8194 370774
rect -7958 370538 -7874 370774
rect -7638 370538 591562 370774
rect 591798 370538 591882 370774
rect 592118 370538 607700 370774
rect -23776 370506 607700 370538
rect -23776 367374 607700 367406
rect -23776 367138 -5084 367374
rect -4848 367138 -4764 367374
rect -4528 367138 7876 367374
rect 8112 367138 8196 367374
rect 8432 367138 38032 367374
rect 38268 367138 38352 367374
rect 38588 367138 74032 367374
rect 74268 367138 74352 367374
rect 74588 367138 110032 367374
rect 110268 367138 110352 367374
rect 110588 367138 146032 367374
rect 146268 367138 146352 367374
rect 146588 367138 182032 367374
rect 182268 367138 182352 367374
rect 182588 367138 218032 367374
rect 218268 367138 218352 367374
rect 218588 367138 254032 367374
rect 254268 367138 254352 367374
rect 254588 367138 290032 367374
rect 290268 367138 290352 367374
rect 290588 367138 326032 367374
rect 326268 367138 326352 367374
rect 326588 367138 362032 367374
rect 362268 367138 362352 367374
rect 362588 367138 398032 367374
rect 398268 367138 398352 367374
rect 398588 367138 434032 367374
rect 434268 367138 434352 367374
rect 434588 367138 470032 367374
rect 470268 367138 470352 367374
rect 470588 367138 506032 367374
rect 506268 367138 506352 367374
rect 506588 367138 542032 367374
rect 542268 367138 542352 367374
rect 542588 367138 571532 367374
rect 571768 367138 571852 367374
rect 572088 367138 588452 367374
rect 588688 367138 588772 367374
rect 589008 367138 607700 367374
rect -23776 367054 607700 367138
rect -23776 366818 -5084 367054
rect -4848 366818 -4764 367054
rect -4528 366818 7876 367054
rect 8112 366818 8196 367054
rect 8432 366818 38032 367054
rect 38268 366818 38352 367054
rect 38588 366818 74032 367054
rect 74268 366818 74352 367054
rect 74588 366818 110032 367054
rect 110268 366818 110352 367054
rect 110588 366818 146032 367054
rect 146268 366818 146352 367054
rect 146588 366818 182032 367054
rect 182268 366818 182352 367054
rect 182588 366818 218032 367054
rect 218268 366818 218352 367054
rect 218588 366818 254032 367054
rect 254268 366818 254352 367054
rect 254588 366818 290032 367054
rect 290268 366818 290352 367054
rect 290588 366818 326032 367054
rect 326268 366818 326352 367054
rect 326588 366818 362032 367054
rect 362268 366818 362352 367054
rect 362588 366818 398032 367054
rect 398268 366818 398352 367054
rect 398588 366818 434032 367054
rect 434268 366818 434352 367054
rect 434588 366818 470032 367054
rect 470268 366818 470352 367054
rect 470588 366818 506032 367054
rect 506268 366818 506352 367054
rect 506588 366818 542032 367054
rect 542268 366818 542352 367054
rect 542588 366818 571532 367054
rect 571768 366818 571852 367054
rect 572088 366818 588452 367054
rect 588688 366818 588772 367054
rect 589008 366818 607700 367054
rect -23776 366786 607700 366818
rect -23776 363654 607700 363686
rect -23776 363418 -1974 363654
rect -1738 363418 -1654 363654
rect -1418 363418 9116 363654
rect 9352 363418 9436 363654
rect 9672 363418 56652 363654
rect 56888 363418 56972 363654
rect 57208 363418 92652 363654
rect 92888 363418 92972 363654
rect 93208 363418 128652 363654
rect 128888 363418 128972 363654
rect 129208 363418 164652 363654
rect 164888 363418 164972 363654
rect 165208 363418 200652 363654
rect 200888 363418 200972 363654
rect 201208 363418 236652 363654
rect 236888 363418 236972 363654
rect 237208 363418 272652 363654
rect 272888 363418 272972 363654
rect 273208 363418 308652 363654
rect 308888 363418 308972 363654
rect 309208 363418 344652 363654
rect 344888 363418 344972 363654
rect 345208 363418 380652 363654
rect 380888 363418 380972 363654
rect 381208 363418 416652 363654
rect 416888 363418 416972 363654
rect 417208 363418 452652 363654
rect 452888 363418 452972 363654
rect 453208 363418 488652 363654
rect 488888 363418 488972 363654
rect 489208 363418 524652 363654
rect 524888 363418 524972 363654
rect 525208 363418 560652 363654
rect 560888 363418 560972 363654
rect 561208 363418 570292 363654
rect 570528 363418 570612 363654
rect 570848 363418 585342 363654
rect 585578 363418 585662 363654
rect 585898 363418 607700 363654
rect -23776 363334 607700 363418
rect -23776 363098 -1974 363334
rect -1738 363098 -1654 363334
rect -1418 363098 9116 363334
rect 9352 363098 9436 363334
rect 9672 363098 56652 363334
rect 56888 363098 56972 363334
rect 57208 363098 92652 363334
rect 92888 363098 92972 363334
rect 93208 363098 128652 363334
rect 128888 363098 128972 363334
rect 129208 363098 164652 363334
rect 164888 363098 164972 363334
rect 165208 363098 200652 363334
rect 200888 363098 200972 363334
rect 201208 363098 236652 363334
rect 236888 363098 236972 363334
rect 237208 363098 272652 363334
rect 272888 363098 272972 363334
rect 273208 363098 308652 363334
rect 308888 363098 308972 363334
rect 309208 363098 344652 363334
rect 344888 363098 344972 363334
rect 345208 363098 380652 363334
rect 380888 363098 380972 363334
rect 381208 363098 416652 363334
rect 416888 363098 416972 363334
rect 417208 363098 452652 363334
rect 452888 363098 452972 363334
rect 453208 363098 488652 363334
rect 488888 363098 488972 363334
rect 489208 363098 524652 363334
rect 524888 363098 524972 363334
rect 525208 363098 560652 363334
rect 560888 363098 560972 363334
rect 561208 363098 570292 363334
rect 570528 363098 570612 363334
rect 570848 363098 585342 363334
rect 585578 363098 585662 363334
rect 585898 363098 607700 363334
rect -23776 363066 607700 363098
rect -23776 349694 607700 349726
rect -23776 349458 -23744 349694
rect -23508 349458 -23424 349694
rect -23188 349458 607112 349694
rect 607348 349458 607432 349694
rect 607668 349458 607700 349694
rect -23776 349374 607700 349458
rect -23776 349138 -23744 349374
rect -23508 349138 -23424 349374
rect -23188 349138 607112 349374
rect 607348 349138 607432 349374
rect 607668 349138 607700 349374
rect -23776 349106 607700 349138
rect -23776 345974 607700 346006
rect -23776 345738 -20634 345974
rect -20398 345738 -20314 345974
rect -20078 345738 604002 345974
rect 604238 345738 604322 345974
rect 604558 345738 607700 345974
rect -23776 345654 607700 345738
rect -23776 345418 -20634 345654
rect -20398 345418 -20314 345654
rect -20078 345418 604002 345654
rect 604238 345418 604322 345654
rect 604558 345418 607700 345654
rect -23776 345386 607700 345418
rect -23776 342254 607700 342286
rect -23776 342018 -17524 342254
rect -17288 342018 -17204 342254
rect -16968 342018 580626 342254
rect 580862 342018 580946 342254
rect 581182 342018 600892 342254
rect 601128 342018 601212 342254
rect 601448 342018 607700 342254
rect -23776 341934 607700 342018
rect -23776 341698 -17524 341934
rect -17288 341698 -17204 341934
rect -16968 341698 580626 341934
rect 580862 341698 580946 341934
rect 581182 341698 600892 341934
rect 601128 341698 601212 341934
rect 601448 341698 607700 341934
rect -23776 341666 607700 341698
rect -23776 338534 607700 338566
rect -23776 338298 -14414 338534
rect -14178 338298 -14094 338534
rect -13858 338298 597782 338534
rect 598018 338298 598102 338534
rect 598338 338298 607700 338534
rect -23776 338214 607700 338298
rect -23776 337978 -14414 338214
rect -14178 337978 -14094 338214
rect -13858 337978 597782 338214
rect 598018 337978 598102 338214
rect 598338 337978 607700 338214
rect -23776 337946 607700 337978
rect -23776 334814 607700 334846
rect -23776 334578 -11304 334814
rect -11068 334578 -10984 334814
rect -10748 334578 594672 334814
rect 594908 334578 594992 334814
rect 595228 334578 607700 334814
rect -23776 334494 607700 334578
rect -23776 334258 -11304 334494
rect -11068 334258 -10984 334494
rect -10748 334258 594672 334494
rect 594908 334258 594992 334494
rect 595228 334258 607700 334494
rect -23776 334226 607700 334258
rect -23776 331094 607700 331126
rect -23776 330858 -8194 331094
rect -7958 330858 -7874 331094
rect -7638 330858 591562 331094
rect 591798 330858 591882 331094
rect 592118 330858 607700 331094
rect -23776 330774 607700 330858
rect -23776 330538 -8194 330774
rect -7958 330538 -7874 330774
rect -7638 330538 591562 330774
rect 591798 330538 591882 330774
rect 592118 330538 607700 330774
rect -23776 330506 607700 330538
rect -23776 327374 607700 327406
rect -23776 327138 -5084 327374
rect -4848 327138 -4764 327374
rect -4528 327138 7876 327374
rect 8112 327138 8196 327374
rect 8432 327138 38032 327374
rect 38268 327138 38352 327374
rect 38588 327138 74032 327374
rect 74268 327138 74352 327374
rect 74588 327138 110032 327374
rect 110268 327138 110352 327374
rect 110588 327138 146032 327374
rect 146268 327138 146352 327374
rect 146588 327138 182032 327374
rect 182268 327138 182352 327374
rect 182588 327138 218032 327374
rect 218268 327138 218352 327374
rect 218588 327138 254032 327374
rect 254268 327138 254352 327374
rect 254588 327138 290032 327374
rect 290268 327138 290352 327374
rect 290588 327138 326032 327374
rect 326268 327138 326352 327374
rect 326588 327138 362032 327374
rect 362268 327138 362352 327374
rect 362588 327138 398032 327374
rect 398268 327138 398352 327374
rect 398588 327138 434032 327374
rect 434268 327138 434352 327374
rect 434588 327138 470032 327374
rect 470268 327138 470352 327374
rect 470588 327138 506032 327374
rect 506268 327138 506352 327374
rect 506588 327138 542032 327374
rect 542268 327138 542352 327374
rect 542588 327138 571532 327374
rect 571768 327138 571852 327374
rect 572088 327138 588452 327374
rect 588688 327138 588772 327374
rect 589008 327138 607700 327374
rect -23776 327054 607700 327138
rect -23776 326818 -5084 327054
rect -4848 326818 -4764 327054
rect -4528 326818 7876 327054
rect 8112 326818 8196 327054
rect 8432 326818 38032 327054
rect 38268 326818 38352 327054
rect 38588 326818 74032 327054
rect 74268 326818 74352 327054
rect 74588 326818 110032 327054
rect 110268 326818 110352 327054
rect 110588 326818 146032 327054
rect 146268 326818 146352 327054
rect 146588 326818 182032 327054
rect 182268 326818 182352 327054
rect 182588 326818 218032 327054
rect 218268 326818 218352 327054
rect 218588 326818 254032 327054
rect 254268 326818 254352 327054
rect 254588 326818 290032 327054
rect 290268 326818 290352 327054
rect 290588 326818 326032 327054
rect 326268 326818 326352 327054
rect 326588 326818 362032 327054
rect 362268 326818 362352 327054
rect 362588 326818 398032 327054
rect 398268 326818 398352 327054
rect 398588 326818 434032 327054
rect 434268 326818 434352 327054
rect 434588 326818 470032 327054
rect 470268 326818 470352 327054
rect 470588 326818 506032 327054
rect 506268 326818 506352 327054
rect 506588 326818 542032 327054
rect 542268 326818 542352 327054
rect 542588 326818 571532 327054
rect 571768 326818 571852 327054
rect 572088 326818 588452 327054
rect 588688 326818 588772 327054
rect 589008 326818 607700 327054
rect -23776 326786 607700 326818
rect -23776 323654 607700 323686
rect -23776 323418 -1974 323654
rect -1738 323418 -1654 323654
rect -1418 323418 9116 323654
rect 9352 323418 9436 323654
rect 9672 323418 56652 323654
rect 56888 323418 56972 323654
rect 57208 323418 92652 323654
rect 92888 323418 92972 323654
rect 93208 323418 128652 323654
rect 128888 323418 128972 323654
rect 129208 323418 164652 323654
rect 164888 323418 164972 323654
rect 165208 323418 200652 323654
rect 200888 323418 200972 323654
rect 201208 323418 236652 323654
rect 236888 323418 236972 323654
rect 237208 323418 272652 323654
rect 272888 323418 272972 323654
rect 273208 323418 308652 323654
rect 308888 323418 308972 323654
rect 309208 323418 344652 323654
rect 344888 323418 344972 323654
rect 345208 323418 380652 323654
rect 380888 323418 380972 323654
rect 381208 323418 416652 323654
rect 416888 323418 416972 323654
rect 417208 323418 452652 323654
rect 452888 323418 452972 323654
rect 453208 323418 488652 323654
rect 488888 323418 488972 323654
rect 489208 323418 524652 323654
rect 524888 323418 524972 323654
rect 525208 323418 560652 323654
rect 560888 323418 560972 323654
rect 561208 323418 570292 323654
rect 570528 323418 570612 323654
rect 570848 323418 585342 323654
rect 585578 323418 585662 323654
rect 585898 323418 607700 323654
rect -23776 323334 607700 323418
rect -23776 323098 -1974 323334
rect -1738 323098 -1654 323334
rect -1418 323098 9116 323334
rect 9352 323098 9436 323334
rect 9672 323098 56652 323334
rect 56888 323098 56972 323334
rect 57208 323098 92652 323334
rect 92888 323098 92972 323334
rect 93208 323098 128652 323334
rect 128888 323098 128972 323334
rect 129208 323098 164652 323334
rect 164888 323098 164972 323334
rect 165208 323098 200652 323334
rect 200888 323098 200972 323334
rect 201208 323098 236652 323334
rect 236888 323098 236972 323334
rect 237208 323098 272652 323334
rect 272888 323098 272972 323334
rect 273208 323098 308652 323334
rect 308888 323098 308972 323334
rect 309208 323098 344652 323334
rect 344888 323098 344972 323334
rect 345208 323098 380652 323334
rect 380888 323098 380972 323334
rect 381208 323098 416652 323334
rect 416888 323098 416972 323334
rect 417208 323098 452652 323334
rect 452888 323098 452972 323334
rect 453208 323098 488652 323334
rect 488888 323098 488972 323334
rect 489208 323098 524652 323334
rect 524888 323098 524972 323334
rect 525208 323098 560652 323334
rect 560888 323098 560972 323334
rect 561208 323098 570292 323334
rect 570528 323098 570612 323334
rect 570848 323098 585342 323334
rect 585578 323098 585662 323334
rect 585898 323098 607700 323334
rect -23776 323066 607700 323098
rect -23776 309694 607700 309726
rect -23776 309458 -23744 309694
rect -23508 309458 -23424 309694
rect -23188 309458 607112 309694
rect 607348 309458 607432 309694
rect 607668 309458 607700 309694
rect -23776 309374 607700 309458
rect -23776 309138 -23744 309374
rect -23508 309138 -23424 309374
rect -23188 309138 607112 309374
rect 607348 309138 607432 309374
rect 607668 309138 607700 309374
rect -23776 309106 607700 309138
rect -23776 305974 607700 306006
rect -23776 305738 -20634 305974
rect -20398 305738 -20314 305974
rect -20078 305738 604002 305974
rect 604238 305738 604322 305974
rect 604558 305738 607700 305974
rect -23776 305654 607700 305738
rect -23776 305418 -20634 305654
rect -20398 305418 -20314 305654
rect -20078 305418 604002 305654
rect 604238 305418 604322 305654
rect 604558 305418 607700 305654
rect -23776 305386 607700 305418
rect -23776 302254 607700 302286
rect -23776 302018 -17524 302254
rect -17288 302018 -17204 302254
rect -16968 302018 580626 302254
rect 580862 302018 580946 302254
rect 581182 302018 600892 302254
rect 601128 302018 601212 302254
rect 601448 302018 607700 302254
rect -23776 301934 607700 302018
rect -23776 301698 -17524 301934
rect -17288 301698 -17204 301934
rect -16968 301698 580626 301934
rect 580862 301698 580946 301934
rect 581182 301698 600892 301934
rect 601128 301698 601212 301934
rect 601448 301698 607700 301934
rect -23776 301666 607700 301698
rect -23776 298534 607700 298566
rect -23776 298298 -14414 298534
rect -14178 298298 -14094 298534
rect -13858 298298 597782 298534
rect 598018 298298 598102 298534
rect 598338 298298 607700 298534
rect -23776 298214 607700 298298
rect -23776 297978 -14414 298214
rect -14178 297978 -14094 298214
rect -13858 297978 597782 298214
rect 598018 297978 598102 298214
rect 598338 297978 607700 298214
rect -23776 297946 607700 297978
rect -23776 294814 607700 294846
rect -23776 294578 -11304 294814
rect -11068 294578 -10984 294814
rect -10748 294578 594672 294814
rect 594908 294578 594992 294814
rect 595228 294578 607700 294814
rect -23776 294494 607700 294578
rect -23776 294258 -11304 294494
rect -11068 294258 -10984 294494
rect -10748 294258 594672 294494
rect 594908 294258 594992 294494
rect 595228 294258 607700 294494
rect -23776 294226 607700 294258
rect -23776 291094 607700 291126
rect -23776 290858 -8194 291094
rect -7958 290858 -7874 291094
rect -7638 290858 591562 291094
rect 591798 290858 591882 291094
rect 592118 290858 607700 291094
rect -23776 290774 607700 290858
rect -23776 290538 -8194 290774
rect -7958 290538 -7874 290774
rect -7638 290538 591562 290774
rect 591798 290538 591882 290774
rect 592118 290538 607700 290774
rect -23776 290506 607700 290538
rect -23776 287374 607700 287406
rect -23776 287138 -5084 287374
rect -4848 287138 -4764 287374
rect -4528 287138 7876 287374
rect 8112 287138 8196 287374
rect 8432 287138 38032 287374
rect 38268 287138 38352 287374
rect 38588 287138 74032 287374
rect 74268 287138 74352 287374
rect 74588 287138 110032 287374
rect 110268 287138 110352 287374
rect 110588 287138 146032 287374
rect 146268 287138 146352 287374
rect 146588 287138 182032 287374
rect 182268 287138 182352 287374
rect 182588 287138 218032 287374
rect 218268 287138 218352 287374
rect 218588 287138 254032 287374
rect 254268 287138 254352 287374
rect 254588 287138 290032 287374
rect 290268 287138 290352 287374
rect 290588 287138 326032 287374
rect 326268 287138 326352 287374
rect 326588 287138 362032 287374
rect 362268 287138 362352 287374
rect 362588 287138 398032 287374
rect 398268 287138 398352 287374
rect 398588 287138 434032 287374
rect 434268 287138 434352 287374
rect 434588 287138 470032 287374
rect 470268 287138 470352 287374
rect 470588 287138 506032 287374
rect 506268 287138 506352 287374
rect 506588 287138 542032 287374
rect 542268 287138 542352 287374
rect 542588 287138 571532 287374
rect 571768 287138 571852 287374
rect 572088 287138 588452 287374
rect 588688 287138 588772 287374
rect 589008 287138 607700 287374
rect -23776 287054 607700 287138
rect -23776 286818 -5084 287054
rect -4848 286818 -4764 287054
rect -4528 286818 7876 287054
rect 8112 286818 8196 287054
rect 8432 286818 38032 287054
rect 38268 286818 38352 287054
rect 38588 286818 74032 287054
rect 74268 286818 74352 287054
rect 74588 286818 110032 287054
rect 110268 286818 110352 287054
rect 110588 286818 146032 287054
rect 146268 286818 146352 287054
rect 146588 286818 182032 287054
rect 182268 286818 182352 287054
rect 182588 286818 218032 287054
rect 218268 286818 218352 287054
rect 218588 286818 254032 287054
rect 254268 286818 254352 287054
rect 254588 286818 290032 287054
rect 290268 286818 290352 287054
rect 290588 286818 326032 287054
rect 326268 286818 326352 287054
rect 326588 286818 362032 287054
rect 362268 286818 362352 287054
rect 362588 286818 398032 287054
rect 398268 286818 398352 287054
rect 398588 286818 434032 287054
rect 434268 286818 434352 287054
rect 434588 286818 470032 287054
rect 470268 286818 470352 287054
rect 470588 286818 506032 287054
rect 506268 286818 506352 287054
rect 506588 286818 542032 287054
rect 542268 286818 542352 287054
rect 542588 286818 571532 287054
rect 571768 286818 571852 287054
rect 572088 286818 588452 287054
rect 588688 286818 588772 287054
rect 589008 286818 607700 287054
rect -23776 286786 607700 286818
rect -23776 283654 607700 283686
rect -23776 283418 -1974 283654
rect -1738 283418 -1654 283654
rect -1418 283418 9116 283654
rect 9352 283418 9436 283654
rect 9672 283418 56652 283654
rect 56888 283418 56972 283654
rect 57208 283418 92652 283654
rect 92888 283418 92972 283654
rect 93208 283418 128652 283654
rect 128888 283418 128972 283654
rect 129208 283418 164652 283654
rect 164888 283418 164972 283654
rect 165208 283418 200652 283654
rect 200888 283418 200972 283654
rect 201208 283418 236652 283654
rect 236888 283418 236972 283654
rect 237208 283418 272652 283654
rect 272888 283418 272972 283654
rect 273208 283418 308652 283654
rect 308888 283418 308972 283654
rect 309208 283418 344652 283654
rect 344888 283418 344972 283654
rect 345208 283418 380652 283654
rect 380888 283418 380972 283654
rect 381208 283418 416652 283654
rect 416888 283418 416972 283654
rect 417208 283418 452652 283654
rect 452888 283418 452972 283654
rect 453208 283418 488652 283654
rect 488888 283418 488972 283654
rect 489208 283418 524652 283654
rect 524888 283418 524972 283654
rect 525208 283418 560652 283654
rect 560888 283418 560972 283654
rect 561208 283418 570292 283654
rect 570528 283418 570612 283654
rect 570848 283418 585342 283654
rect 585578 283418 585662 283654
rect 585898 283418 607700 283654
rect -23776 283334 607700 283418
rect -23776 283098 -1974 283334
rect -1738 283098 -1654 283334
rect -1418 283098 9116 283334
rect 9352 283098 9436 283334
rect 9672 283098 56652 283334
rect 56888 283098 56972 283334
rect 57208 283098 92652 283334
rect 92888 283098 92972 283334
rect 93208 283098 128652 283334
rect 128888 283098 128972 283334
rect 129208 283098 164652 283334
rect 164888 283098 164972 283334
rect 165208 283098 200652 283334
rect 200888 283098 200972 283334
rect 201208 283098 236652 283334
rect 236888 283098 236972 283334
rect 237208 283098 272652 283334
rect 272888 283098 272972 283334
rect 273208 283098 308652 283334
rect 308888 283098 308972 283334
rect 309208 283098 344652 283334
rect 344888 283098 344972 283334
rect 345208 283098 380652 283334
rect 380888 283098 380972 283334
rect 381208 283098 416652 283334
rect 416888 283098 416972 283334
rect 417208 283098 452652 283334
rect 452888 283098 452972 283334
rect 453208 283098 488652 283334
rect 488888 283098 488972 283334
rect 489208 283098 524652 283334
rect 524888 283098 524972 283334
rect 525208 283098 560652 283334
rect 560888 283098 560972 283334
rect 561208 283098 570292 283334
rect 570528 283098 570612 283334
rect 570848 283098 585342 283334
rect 585578 283098 585662 283334
rect 585898 283098 607700 283334
rect -23776 283066 607700 283098
rect -23776 269694 607700 269726
rect -23776 269458 -23744 269694
rect -23508 269458 -23424 269694
rect -23188 269458 607112 269694
rect 607348 269458 607432 269694
rect 607668 269458 607700 269694
rect -23776 269374 607700 269458
rect -23776 269138 -23744 269374
rect -23508 269138 -23424 269374
rect -23188 269138 607112 269374
rect 607348 269138 607432 269374
rect 607668 269138 607700 269374
rect -23776 269106 607700 269138
rect -23776 265974 607700 266006
rect -23776 265738 -20634 265974
rect -20398 265738 -20314 265974
rect -20078 265738 604002 265974
rect 604238 265738 604322 265974
rect 604558 265738 607700 265974
rect -23776 265654 607700 265738
rect -23776 265418 -20634 265654
rect -20398 265418 -20314 265654
rect -20078 265418 604002 265654
rect 604238 265418 604322 265654
rect 604558 265418 607700 265654
rect -23776 265386 607700 265418
rect -23776 262254 607700 262286
rect -23776 262018 -17524 262254
rect -17288 262018 -17204 262254
rect -16968 262018 580626 262254
rect 580862 262018 580946 262254
rect 581182 262018 600892 262254
rect 601128 262018 601212 262254
rect 601448 262018 607700 262254
rect -23776 261934 607700 262018
rect -23776 261698 -17524 261934
rect -17288 261698 -17204 261934
rect -16968 261698 580626 261934
rect 580862 261698 580946 261934
rect 581182 261698 600892 261934
rect 601128 261698 601212 261934
rect 601448 261698 607700 261934
rect -23776 261666 607700 261698
rect -23776 258534 607700 258566
rect -23776 258298 -14414 258534
rect -14178 258298 -14094 258534
rect -13858 258298 597782 258534
rect 598018 258298 598102 258534
rect 598338 258298 607700 258534
rect -23776 258214 607700 258298
rect -23776 257978 -14414 258214
rect -14178 257978 -14094 258214
rect -13858 257978 597782 258214
rect 598018 257978 598102 258214
rect 598338 257978 607700 258214
rect -23776 257946 607700 257978
rect -23776 254814 607700 254846
rect -23776 254578 -11304 254814
rect -11068 254578 -10984 254814
rect -10748 254578 594672 254814
rect 594908 254578 594992 254814
rect 595228 254578 607700 254814
rect -23776 254494 607700 254578
rect -23776 254258 -11304 254494
rect -11068 254258 -10984 254494
rect -10748 254258 594672 254494
rect 594908 254258 594992 254494
rect 595228 254258 607700 254494
rect -23776 254226 607700 254258
rect -23776 251094 607700 251126
rect -23776 250858 -8194 251094
rect -7958 250858 -7874 251094
rect -7638 250858 591562 251094
rect 591798 250858 591882 251094
rect 592118 250858 607700 251094
rect -23776 250774 607700 250858
rect -23776 250538 -8194 250774
rect -7958 250538 -7874 250774
rect -7638 250538 591562 250774
rect 591798 250538 591882 250774
rect 592118 250538 607700 250774
rect -23776 250506 607700 250538
rect -23776 247374 607700 247406
rect -23776 247138 -5084 247374
rect -4848 247138 -4764 247374
rect -4528 247138 7876 247374
rect 8112 247138 8196 247374
rect 8432 247138 38032 247374
rect 38268 247138 38352 247374
rect 38588 247138 74032 247374
rect 74268 247138 74352 247374
rect 74588 247138 110032 247374
rect 110268 247138 110352 247374
rect 110588 247138 146032 247374
rect 146268 247138 146352 247374
rect 146588 247138 182032 247374
rect 182268 247138 182352 247374
rect 182588 247138 218032 247374
rect 218268 247138 218352 247374
rect 218588 247138 254032 247374
rect 254268 247138 254352 247374
rect 254588 247138 290032 247374
rect 290268 247138 290352 247374
rect 290588 247138 326032 247374
rect 326268 247138 326352 247374
rect 326588 247138 362032 247374
rect 362268 247138 362352 247374
rect 362588 247138 398032 247374
rect 398268 247138 398352 247374
rect 398588 247138 434032 247374
rect 434268 247138 434352 247374
rect 434588 247138 470032 247374
rect 470268 247138 470352 247374
rect 470588 247138 506032 247374
rect 506268 247138 506352 247374
rect 506588 247138 542032 247374
rect 542268 247138 542352 247374
rect 542588 247138 571532 247374
rect 571768 247138 571852 247374
rect 572088 247138 588452 247374
rect 588688 247138 588772 247374
rect 589008 247138 607700 247374
rect -23776 247054 607700 247138
rect -23776 246818 -5084 247054
rect -4848 246818 -4764 247054
rect -4528 246818 7876 247054
rect 8112 246818 8196 247054
rect 8432 246818 38032 247054
rect 38268 246818 38352 247054
rect 38588 246818 74032 247054
rect 74268 246818 74352 247054
rect 74588 246818 110032 247054
rect 110268 246818 110352 247054
rect 110588 246818 146032 247054
rect 146268 246818 146352 247054
rect 146588 246818 182032 247054
rect 182268 246818 182352 247054
rect 182588 246818 218032 247054
rect 218268 246818 218352 247054
rect 218588 246818 254032 247054
rect 254268 246818 254352 247054
rect 254588 246818 290032 247054
rect 290268 246818 290352 247054
rect 290588 246818 326032 247054
rect 326268 246818 326352 247054
rect 326588 246818 362032 247054
rect 362268 246818 362352 247054
rect 362588 246818 398032 247054
rect 398268 246818 398352 247054
rect 398588 246818 434032 247054
rect 434268 246818 434352 247054
rect 434588 246818 470032 247054
rect 470268 246818 470352 247054
rect 470588 246818 506032 247054
rect 506268 246818 506352 247054
rect 506588 246818 542032 247054
rect 542268 246818 542352 247054
rect 542588 246818 571532 247054
rect 571768 246818 571852 247054
rect 572088 246818 588452 247054
rect 588688 246818 588772 247054
rect 589008 246818 607700 247054
rect -23776 246786 607700 246818
rect -23776 243654 607700 243686
rect -23776 243418 -1974 243654
rect -1738 243418 -1654 243654
rect -1418 243418 9116 243654
rect 9352 243418 9436 243654
rect 9672 243418 56652 243654
rect 56888 243418 56972 243654
rect 57208 243418 92652 243654
rect 92888 243418 92972 243654
rect 93208 243418 128652 243654
rect 128888 243418 128972 243654
rect 129208 243418 164652 243654
rect 164888 243418 164972 243654
rect 165208 243418 200652 243654
rect 200888 243418 200972 243654
rect 201208 243418 236652 243654
rect 236888 243418 236972 243654
rect 237208 243418 272652 243654
rect 272888 243418 272972 243654
rect 273208 243418 308652 243654
rect 308888 243418 308972 243654
rect 309208 243418 344652 243654
rect 344888 243418 344972 243654
rect 345208 243418 380652 243654
rect 380888 243418 380972 243654
rect 381208 243418 416652 243654
rect 416888 243418 416972 243654
rect 417208 243418 452652 243654
rect 452888 243418 452972 243654
rect 453208 243418 488652 243654
rect 488888 243418 488972 243654
rect 489208 243418 524652 243654
rect 524888 243418 524972 243654
rect 525208 243418 560652 243654
rect 560888 243418 560972 243654
rect 561208 243418 570292 243654
rect 570528 243418 570612 243654
rect 570848 243418 585342 243654
rect 585578 243418 585662 243654
rect 585898 243418 607700 243654
rect -23776 243334 607700 243418
rect -23776 243098 -1974 243334
rect -1738 243098 -1654 243334
rect -1418 243098 9116 243334
rect 9352 243098 9436 243334
rect 9672 243098 56652 243334
rect 56888 243098 56972 243334
rect 57208 243098 92652 243334
rect 92888 243098 92972 243334
rect 93208 243098 128652 243334
rect 128888 243098 128972 243334
rect 129208 243098 164652 243334
rect 164888 243098 164972 243334
rect 165208 243098 200652 243334
rect 200888 243098 200972 243334
rect 201208 243098 236652 243334
rect 236888 243098 236972 243334
rect 237208 243098 272652 243334
rect 272888 243098 272972 243334
rect 273208 243098 308652 243334
rect 308888 243098 308972 243334
rect 309208 243098 344652 243334
rect 344888 243098 344972 243334
rect 345208 243098 380652 243334
rect 380888 243098 380972 243334
rect 381208 243098 416652 243334
rect 416888 243098 416972 243334
rect 417208 243098 452652 243334
rect 452888 243098 452972 243334
rect 453208 243098 488652 243334
rect 488888 243098 488972 243334
rect 489208 243098 524652 243334
rect 524888 243098 524972 243334
rect 525208 243098 560652 243334
rect 560888 243098 560972 243334
rect 561208 243098 570292 243334
rect 570528 243098 570612 243334
rect 570848 243098 585342 243334
rect 585578 243098 585662 243334
rect 585898 243098 607700 243334
rect -23776 243066 607700 243098
rect -23776 229694 607700 229726
rect -23776 229458 -23744 229694
rect -23508 229458 -23424 229694
rect -23188 229458 607112 229694
rect 607348 229458 607432 229694
rect 607668 229458 607700 229694
rect -23776 229374 607700 229458
rect -23776 229138 -23744 229374
rect -23508 229138 -23424 229374
rect -23188 229138 607112 229374
rect 607348 229138 607432 229374
rect 607668 229138 607700 229374
rect -23776 229106 607700 229138
rect -23776 225974 607700 226006
rect -23776 225738 -20634 225974
rect -20398 225738 -20314 225974
rect -20078 225738 604002 225974
rect 604238 225738 604322 225974
rect 604558 225738 607700 225974
rect -23776 225654 607700 225738
rect -23776 225418 -20634 225654
rect -20398 225418 -20314 225654
rect -20078 225418 604002 225654
rect 604238 225418 604322 225654
rect 604558 225418 607700 225654
rect -23776 225386 607700 225418
rect -23776 222254 607700 222286
rect -23776 222018 -17524 222254
rect -17288 222018 -17204 222254
rect -16968 222018 580626 222254
rect 580862 222018 580946 222254
rect 581182 222018 600892 222254
rect 601128 222018 601212 222254
rect 601448 222018 607700 222254
rect -23776 221934 607700 222018
rect -23776 221698 -17524 221934
rect -17288 221698 -17204 221934
rect -16968 221698 580626 221934
rect 580862 221698 580946 221934
rect 581182 221698 600892 221934
rect 601128 221698 601212 221934
rect 601448 221698 607700 221934
rect -23776 221666 607700 221698
rect -23776 218534 607700 218566
rect -23776 218298 -14414 218534
rect -14178 218298 -14094 218534
rect -13858 218298 597782 218534
rect 598018 218298 598102 218534
rect 598338 218298 607700 218534
rect -23776 218214 607700 218298
rect -23776 217978 -14414 218214
rect -14178 217978 -14094 218214
rect -13858 217978 597782 218214
rect 598018 217978 598102 218214
rect 598338 217978 607700 218214
rect -23776 217946 607700 217978
rect -23776 214814 607700 214846
rect -23776 214578 -11304 214814
rect -11068 214578 -10984 214814
rect -10748 214578 594672 214814
rect 594908 214578 594992 214814
rect 595228 214578 607700 214814
rect -23776 214494 607700 214578
rect -23776 214258 -11304 214494
rect -11068 214258 -10984 214494
rect -10748 214258 594672 214494
rect 594908 214258 594992 214494
rect 595228 214258 607700 214494
rect -23776 214226 607700 214258
rect -23776 211094 607700 211126
rect -23776 210858 -8194 211094
rect -7958 210858 -7874 211094
rect -7638 210858 591562 211094
rect 591798 210858 591882 211094
rect 592118 210858 607700 211094
rect -23776 210774 607700 210858
rect -23776 210538 -8194 210774
rect -7958 210538 -7874 210774
rect -7638 210538 591562 210774
rect 591798 210538 591882 210774
rect 592118 210538 607700 210774
rect -23776 210506 607700 210538
rect -23776 207374 607700 207406
rect -23776 207138 -5084 207374
rect -4848 207138 -4764 207374
rect -4528 207138 7876 207374
rect 8112 207138 8196 207374
rect 8432 207138 38032 207374
rect 38268 207138 38352 207374
rect 38588 207138 74032 207374
rect 74268 207138 74352 207374
rect 74588 207138 110032 207374
rect 110268 207138 110352 207374
rect 110588 207138 146032 207374
rect 146268 207138 146352 207374
rect 146588 207138 182032 207374
rect 182268 207138 182352 207374
rect 182588 207138 218032 207374
rect 218268 207138 218352 207374
rect 218588 207138 254032 207374
rect 254268 207138 254352 207374
rect 254588 207138 290032 207374
rect 290268 207138 290352 207374
rect 290588 207138 326032 207374
rect 326268 207138 326352 207374
rect 326588 207138 362032 207374
rect 362268 207138 362352 207374
rect 362588 207138 398032 207374
rect 398268 207138 398352 207374
rect 398588 207138 434032 207374
rect 434268 207138 434352 207374
rect 434588 207138 470032 207374
rect 470268 207138 470352 207374
rect 470588 207138 506032 207374
rect 506268 207138 506352 207374
rect 506588 207138 542032 207374
rect 542268 207138 542352 207374
rect 542588 207138 571532 207374
rect 571768 207138 571852 207374
rect 572088 207138 588452 207374
rect 588688 207138 588772 207374
rect 589008 207138 607700 207374
rect -23776 207054 607700 207138
rect -23776 206818 -5084 207054
rect -4848 206818 -4764 207054
rect -4528 206818 7876 207054
rect 8112 206818 8196 207054
rect 8432 206818 38032 207054
rect 38268 206818 38352 207054
rect 38588 206818 74032 207054
rect 74268 206818 74352 207054
rect 74588 206818 110032 207054
rect 110268 206818 110352 207054
rect 110588 206818 146032 207054
rect 146268 206818 146352 207054
rect 146588 206818 182032 207054
rect 182268 206818 182352 207054
rect 182588 206818 218032 207054
rect 218268 206818 218352 207054
rect 218588 206818 254032 207054
rect 254268 206818 254352 207054
rect 254588 206818 290032 207054
rect 290268 206818 290352 207054
rect 290588 206818 326032 207054
rect 326268 206818 326352 207054
rect 326588 206818 362032 207054
rect 362268 206818 362352 207054
rect 362588 206818 398032 207054
rect 398268 206818 398352 207054
rect 398588 206818 434032 207054
rect 434268 206818 434352 207054
rect 434588 206818 470032 207054
rect 470268 206818 470352 207054
rect 470588 206818 506032 207054
rect 506268 206818 506352 207054
rect 506588 206818 542032 207054
rect 542268 206818 542352 207054
rect 542588 206818 571532 207054
rect 571768 206818 571852 207054
rect 572088 206818 588452 207054
rect 588688 206818 588772 207054
rect 589008 206818 607700 207054
rect -23776 206786 607700 206818
rect -23776 203654 607700 203686
rect -23776 203418 -1974 203654
rect -1738 203418 -1654 203654
rect -1418 203418 9116 203654
rect 9352 203418 9436 203654
rect 9672 203418 56652 203654
rect 56888 203418 56972 203654
rect 57208 203418 92652 203654
rect 92888 203418 92972 203654
rect 93208 203418 128652 203654
rect 128888 203418 128972 203654
rect 129208 203418 164652 203654
rect 164888 203418 164972 203654
rect 165208 203418 200652 203654
rect 200888 203418 200972 203654
rect 201208 203418 236652 203654
rect 236888 203418 236972 203654
rect 237208 203418 272652 203654
rect 272888 203418 272972 203654
rect 273208 203418 308652 203654
rect 308888 203418 308972 203654
rect 309208 203418 344652 203654
rect 344888 203418 344972 203654
rect 345208 203418 380652 203654
rect 380888 203418 380972 203654
rect 381208 203418 416652 203654
rect 416888 203418 416972 203654
rect 417208 203418 452652 203654
rect 452888 203418 452972 203654
rect 453208 203418 488652 203654
rect 488888 203418 488972 203654
rect 489208 203418 524652 203654
rect 524888 203418 524972 203654
rect 525208 203418 560652 203654
rect 560888 203418 560972 203654
rect 561208 203418 570292 203654
rect 570528 203418 570612 203654
rect 570848 203418 585342 203654
rect 585578 203418 585662 203654
rect 585898 203418 607700 203654
rect -23776 203334 607700 203418
rect -23776 203098 -1974 203334
rect -1738 203098 -1654 203334
rect -1418 203098 9116 203334
rect 9352 203098 9436 203334
rect 9672 203098 56652 203334
rect 56888 203098 56972 203334
rect 57208 203098 92652 203334
rect 92888 203098 92972 203334
rect 93208 203098 128652 203334
rect 128888 203098 128972 203334
rect 129208 203098 164652 203334
rect 164888 203098 164972 203334
rect 165208 203098 200652 203334
rect 200888 203098 200972 203334
rect 201208 203098 236652 203334
rect 236888 203098 236972 203334
rect 237208 203098 272652 203334
rect 272888 203098 272972 203334
rect 273208 203098 308652 203334
rect 308888 203098 308972 203334
rect 309208 203098 344652 203334
rect 344888 203098 344972 203334
rect 345208 203098 380652 203334
rect 380888 203098 380972 203334
rect 381208 203098 416652 203334
rect 416888 203098 416972 203334
rect 417208 203098 452652 203334
rect 452888 203098 452972 203334
rect 453208 203098 488652 203334
rect 488888 203098 488972 203334
rect 489208 203098 524652 203334
rect 524888 203098 524972 203334
rect 525208 203098 560652 203334
rect 560888 203098 560972 203334
rect 561208 203098 570292 203334
rect 570528 203098 570612 203334
rect 570848 203098 585342 203334
rect 585578 203098 585662 203334
rect 585898 203098 607700 203334
rect -23776 203066 607700 203098
rect -23776 189694 607700 189726
rect -23776 189458 -23744 189694
rect -23508 189458 -23424 189694
rect -23188 189458 607112 189694
rect 607348 189458 607432 189694
rect 607668 189458 607700 189694
rect -23776 189374 607700 189458
rect -23776 189138 -23744 189374
rect -23508 189138 -23424 189374
rect -23188 189138 607112 189374
rect 607348 189138 607432 189374
rect 607668 189138 607700 189374
rect -23776 189106 607700 189138
rect -23776 185974 607700 186006
rect -23776 185738 -20634 185974
rect -20398 185738 -20314 185974
rect -20078 185738 604002 185974
rect 604238 185738 604322 185974
rect 604558 185738 607700 185974
rect -23776 185654 607700 185738
rect -23776 185418 -20634 185654
rect -20398 185418 -20314 185654
rect -20078 185418 604002 185654
rect 604238 185418 604322 185654
rect 604558 185418 607700 185654
rect -23776 185386 607700 185418
rect -23776 182254 607700 182286
rect -23776 182018 -17524 182254
rect -17288 182018 -17204 182254
rect -16968 182018 580626 182254
rect 580862 182018 580946 182254
rect 581182 182018 600892 182254
rect 601128 182018 601212 182254
rect 601448 182018 607700 182254
rect -23776 181934 607700 182018
rect -23776 181698 -17524 181934
rect -17288 181698 -17204 181934
rect -16968 181698 580626 181934
rect 580862 181698 580946 181934
rect 581182 181698 600892 181934
rect 601128 181698 601212 181934
rect 601448 181698 607700 181934
rect -23776 181666 607700 181698
rect -23776 178534 607700 178566
rect -23776 178298 -14414 178534
rect -14178 178298 -14094 178534
rect -13858 178298 597782 178534
rect 598018 178298 598102 178534
rect 598338 178298 607700 178534
rect -23776 178214 607700 178298
rect -23776 177978 -14414 178214
rect -14178 177978 -14094 178214
rect -13858 177978 597782 178214
rect 598018 177978 598102 178214
rect 598338 177978 607700 178214
rect -23776 177946 607700 177978
rect -23776 174814 607700 174846
rect -23776 174578 -11304 174814
rect -11068 174578 -10984 174814
rect -10748 174578 594672 174814
rect 594908 174578 594992 174814
rect 595228 174578 607700 174814
rect -23776 174494 607700 174578
rect -23776 174258 -11304 174494
rect -11068 174258 -10984 174494
rect -10748 174258 594672 174494
rect 594908 174258 594992 174494
rect 595228 174258 607700 174494
rect -23776 174226 607700 174258
rect -23776 171094 607700 171126
rect -23776 170858 -8194 171094
rect -7958 170858 -7874 171094
rect -7638 170858 591562 171094
rect 591798 170858 591882 171094
rect 592118 170858 607700 171094
rect -23776 170774 607700 170858
rect -23776 170538 -8194 170774
rect -7958 170538 -7874 170774
rect -7638 170538 591562 170774
rect 591798 170538 591882 170774
rect 592118 170538 607700 170774
rect -23776 170506 607700 170538
rect -23776 167374 607700 167406
rect -23776 167138 -5084 167374
rect -4848 167138 -4764 167374
rect -4528 167138 7876 167374
rect 8112 167138 8196 167374
rect 8432 167138 38032 167374
rect 38268 167138 38352 167374
rect 38588 167138 60622 167374
rect 60858 167138 159098 167374
rect 159334 167138 182032 167374
rect 182268 167138 182352 167374
rect 182588 167138 185622 167374
rect 185858 167138 284098 167374
rect 284334 167138 290032 167374
rect 290268 167138 290352 167374
rect 290588 167138 310622 167374
rect 310858 167138 409098 167374
rect 409334 167138 434032 167374
rect 434268 167138 434352 167374
rect 434588 167138 436622 167374
rect 436858 167138 535098 167374
rect 535334 167138 542032 167374
rect 542268 167138 542352 167374
rect 542588 167138 571532 167374
rect 571768 167138 571852 167374
rect 572088 167138 588452 167374
rect 588688 167138 588772 167374
rect 589008 167138 607700 167374
rect -23776 167054 607700 167138
rect -23776 166818 -5084 167054
rect -4848 166818 -4764 167054
rect -4528 166818 7876 167054
rect 8112 166818 8196 167054
rect 8432 166818 38032 167054
rect 38268 166818 38352 167054
rect 38588 166818 60622 167054
rect 60858 166818 159098 167054
rect 159334 166818 182032 167054
rect 182268 166818 182352 167054
rect 182588 166818 185622 167054
rect 185858 166818 284098 167054
rect 284334 166818 290032 167054
rect 290268 166818 290352 167054
rect 290588 166818 310622 167054
rect 310858 166818 409098 167054
rect 409334 166818 434032 167054
rect 434268 166818 434352 167054
rect 434588 166818 436622 167054
rect 436858 166818 535098 167054
rect 535334 166818 542032 167054
rect 542268 166818 542352 167054
rect 542588 166818 571532 167054
rect 571768 166818 571852 167054
rect 572088 166818 588452 167054
rect 588688 166818 588772 167054
rect 589008 166818 607700 167054
rect -23776 166786 607700 166818
rect -23776 163654 607700 163686
rect -23776 163418 -1974 163654
rect -1738 163418 -1654 163654
rect -1418 163418 9116 163654
rect 9352 163418 9436 163654
rect 9672 163418 56652 163654
rect 56888 163418 56972 163654
rect 57208 163418 61342 163654
rect 61578 163418 158378 163654
rect 158614 163418 164652 163654
rect 164888 163418 164972 163654
rect 165208 163418 186342 163654
rect 186578 163418 283378 163654
rect 283614 163418 308652 163654
rect 308888 163418 308972 163654
rect 309208 163418 311342 163654
rect 311578 163418 408378 163654
rect 408614 163418 416652 163654
rect 416888 163418 416972 163654
rect 417208 163418 437342 163654
rect 437578 163418 534378 163654
rect 534614 163418 560652 163654
rect 560888 163418 560972 163654
rect 561208 163418 570292 163654
rect 570528 163418 570612 163654
rect 570848 163418 585342 163654
rect 585578 163418 585662 163654
rect 585898 163418 607700 163654
rect -23776 163334 607700 163418
rect -23776 163098 -1974 163334
rect -1738 163098 -1654 163334
rect -1418 163098 9116 163334
rect 9352 163098 9436 163334
rect 9672 163098 56652 163334
rect 56888 163098 56972 163334
rect 57208 163098 61342 163334
rect 61578 163098 158378 163334
rect 158614 163098 164652 163334
rect 164888 163098 164972 163334
rect 165208 163098 186342 163334
rect 186578 163098 283378 163334
rect 283614 163098 308652 163334
rect 308888 163098 308972 163334
rect 309208 163098 311342 163334
rect 311578 163098 408378 163334
rect 408614 163098 416652 163334
rect 416888 163098 416972 163334
rect 417208 163098 437342 163334
rect 437578 163098 534378 163334
rect 534614 163098 560652 163334
rect 560888 163098 560972 163334
rect 561208 163098 570292 163334
rect 570528 163098 570612 163334
rect 570848 163098 585342 163334
rect 585578 163098 585662 163334
rect 585898 163098 607700 163334
rect -23776 163066 607700 163098
rect -23776 149694 607700 149726
rect -23776 149458 -23744 149694
rect -23508 149458 -23424 149694
rect -23188 149458 607112 149694
rect 607348 149458 607432 149694
rect 607668 149458 607700 149694
rect -23776 149374 607700 149458
rect -23776 149138 -23744 149374
rect -23508 149138 -23424 149374
rect -23188 149138 607112 149374
rect 607348 149138 607432 149374
rect 607668 149138 607700 149374
rect -23776 149106 607700 149138
rect -23776 145974 607700 146006
rect -23776 145738 -20634 145974
rect -20398 145738 -20314 145974
rect -20078 145738 604002 145974
rect 604238 145738 604322 145974
rect 604558 145738 607700 145974
rect -23776 145654 607700 145738
rect -23776 145418 -20634 145654
rect -20398 145418 -20314 145654
rect -20078 145418 604002 145654
rect 604238 145418 604322 145654
rect 604558 145418 607700 145654
rect -23776 145386 607700 145418
rect -23776 142254 607700 142286
rect -23776 142018 -17524 142254
rect -17288 142018 -17204 142254
rect -16968 142018 580626 142254
rect 580862 142018 580946 142254
rect 581182 142018 600892 142254
rect 601128 142018 601212 142254
rect 601448 142018 607700 142254
rect -23776 141934 607700 142018
rect -23776 141698 -17524 141934
rect -17288 141698 -17204 141934
rect -16968 141698 580626 141934
rect 580862 141698 580946 141934
rect 581182 141698 600892 141934
rect 601128 141698 601212 141934
rect 601448 141698 607700 141934
rect -23776 141666 607700 141698
rect -23776 138534 607700 138566
rect -23776 138298 -14414 138534
rect -14178 138298 -14094 138534
rect -13858 138298 597782 138534
rect 598018 138298 598102 138534
rect 598338 138298 607700 138534
rect -23776 138214 607700 138298
rect -23776 137978 -14414 138214
rect -14178 137978 -14094 138214
rect -13858 137978 597782 138214
rect 598018 137978 598102 138214
rect 598338 137978 607700 138214
rect -23776 137946 607700 137978
rect -23776 134814 607700 134846
rect -23776 134578 -11304 134814
rect -11068 134578 -10984 134814
rect -10748 134578 594672 134814
rect 594908 134578 594992 134814
rect 595228 134578 607700 134814
rect -23776 134494 607700 134578
rect -23776 134258 -11304 134494
rect -11068 134258 -10984 134494
rect -10748 134258 594672 134494
rect 594908 134258 594992 134494
rect 595228 134258 607700 134494
rect -23776 134226 607700 134258
rect -23776 131094 607700 131126
rect -23776 130858 -8194 131094
rect -7958 130858 -7874 131094
rect -7638 130858 591562 131094
rect 591798 130858 591882 131094
rect 592118 130858 607700 131094
rect -23776 130774 607700 130858
rect -23776 130538 -8194 130774
rect -7958 130538 -7874 130774
rect -7638 130538 591562 130774
rect 591798 130538 591882 130774
rect 592118 130538 607700 130774
rect -23776 130506 607700 130538
rect -23776 127374 607700 127406
rect -23776 127138 -5084 127374
rect -4848 127138 -4764 127374
rect -4528 127138 7876 127374
rect 8112 127138 8196 127374
rect 8432 127138 38032 127374
rect 38268 127138 38352 127374
rect 38588 127138 60622 127374
rect 60858 127138 159098 127374
rect 159334 127138 182032 127374
rect 182268 127138 182352 127374
rect 182588 127138 185622 127374
rect 185858 127138 284098 127374
rect 284334 127138 290032 127374
rect 290268 127138 290352 127374
rect 290588 127138 310622 127374
rect 310858 127138 409098 127374
rect 409334 127138 434032 127374
rect 434268 127138 434352 127374
rect 434588 127138 436622 127374
rect 436858 127138 535098 127374
rect 535334 127138 542032 127374
rect 542268 127138 542352 127374
rect 542588 127138 571532 127374
rect 571768 127138 571852 127374
rect 572088 127138 588452 127374
rect 588688 127138 588772 127374
rect 589008 127138 607700 127374
rect -23776 127054 607700 127138
rect -23776 126818 -5084 127054
rect -4848 126818 -4764 127054
rect -4528 126818 7876 127054
rect 8112 126818 8196 127054
rect 8432 126818 38032 127054
rect 38268 126818 38352 127054
rect 38588 126818 60622 127054
rect 60858 126818 159098 127054
rect 159334 126818 182032 127054
rect 182268 126818 182352 127054
rect 182588 126818 185622 127054
rect 185858 126818 284098 127054
rect 284334 126818 290032 127054
rect 290268 126818 290352 127054
rect 290588 126818 310622 127054
rect 310858 126818 409098 127054
rect 409334 126818 434032 127054
rect 434268 126818 434352 127054
rect 434588 126818 436622 127054
rect 436858 126818 535098 127054
rect 535334 126818 542032 127054
rect 542268 126818 542352 127054
rect 542588 126818 571532 127054
rect 571768 126818 571852 127054
rect 572088 126818 588452 127054
rect 588688 126818 588772 127054
rect 589008 126818 607700 127054
rect -23776 126786 607700 126818
rect -23776 123654 607700 123686
rect -23776 123418 -1974 123654
rect -1738 123418 -1654 123654
rect -1418 123418 9116 123654
rect 9352 123418 9436 123654
rect 9672 123418 56652 123654
rect 56888 123418 56972 123654
rect 57208 123418 61342 123654
rect 61578 123418 158378 123654
rect 158614 123418 164652 123654
rect 164888 123418 164972 123654
rect 165208 123418 186342 123654
rect 186578 123418 283378 123654
rect 283614 123418 308652 123654
rect 308888 123418 308972 123654
rect 309208 123418 311342 123654
rect 311578 123418 408378 123654
rect 408614 123418 416652 123654
rect 416888 123418 416972 123654
rect 417208 123418 437342 123654
rect 437578 123418 534378 123654
rect 534614 123418 560652 123654
rect 560888 123418 560972 123654
rect 561208 123418 570292 123654
rect 570528 123418 570612 123654
rect 570848 123418 585342 123654
rect 585578 123418 585662 123654
rect 585898 123418 607700 123654
rect -23776 123334 607700 123418
rect -23776 123098 -1974 123334
rect -1738 123098 -1654 123334
rect -1418 123098 9116 123334
rect 9352 123098 9436 123334
rect 9672 123098 56652 123334
rect 56888 123098 56972 123334
rect 57208 123098 61342 123334
rect 61578 123098 158378 123334
rect 158614 123098 164652 123334
rect 164888 123098 164972 123334
rect 165208 123098 186342 123334
rect 186578 123098 283378 123334
rect 283614 123098 308652 123334
rect 308888 123098 308972 123334
rect 309208 123098 311342 123334
rect 311578 123098 408378 123334
rect 408614 123098 416652 123334
rect 416888 123098 416972 123334
rect 417208 123098 437342 123334
rect 437578 123098 534378 123334
rect 534614 123098 560652 123334
rect 560888 123098 560972 123334
rect 561208 123098 570292 123334
rect 570528 123098 570612 123334
rect 570848 123098 585342 123334
rect 585578 123098 585662 123334
rect 585898 123098 607700 123334
rect -23776 123066 607700 123098
rect 61280 121244 61640 121300
rect 61280 121008 61342 121244
rect 61578 121008 61640 121244
rect 61280 120952 61640 121008
rect 62952 121244 63300 121300
rect 62952 121008 63008 121244
rect 63244 121008 63300 121244
rect 62952 120952 63300 121008
rect 281656 121244 282004 121300
rect 281656 121008 281712 121244
rect 281948 121008 282004 121244
rect 281656 120952 282004 121008
rect 283316 121244 283676 121300
rect 283316 121008 283378 121244
rect 283614 121008 283676 121244
rect 283316 120952 283676 121008
rect 311280 121244 311640 121300
rect 311280 121008 311342 121244
rect 311578 121008 311640 121244
rect 311280 120952 311640 121008
rect 312952 121244 313300 121300
rect 312952 121008 313008 121244
rect 313244 121008 313300 121244
rect 312952 120952 313300 121008
rect 532656 121244 533004 121300
rect 532656 121008 532712 121244
rect 532948 121008 533004 121244
rect 532656 120952 533004 121008
rect 534316 121244 534676 121300
rect 534316 121008 534378 121244
rect 534614 121008 534676 121244
rect 534316 120952 534676 121008
rect 157336 120564 157684 120620
rect 157336 120328 157392 120564
rect 157628 120328 157684 120564
rect 157336 120272 157684 120328
rect 159036 120564 159396 120620
rect 159036 120328 159098 120564
rect 159334 120328 159396 120564
rect 159036 120272 159396 120328
rect 185560 120564 185920 120620
rect 185560 120328 185622 120564
rect 185858 120328 185920 120564
rect 185560 120272 185920 120328
rect 187272 120564 187620 120620
rect 187272 120328 187328 120564
rect 187564 120328 187620 120564
rect 187272 120272 187620 120328
rect 407336 120564 407684 120620
rect 407336 120328 407392 120564
rect 407628 120328 407684 120564
rect 407336 120272 407684 120328
rect 409036 120564 409396 120620
rect 409036 120328 409098 120564
rect 409334 120328 409396 120564
rect 409036 120272 409396 120328
rect 436560 120564 436920 120620
rect 436560 120328 436622 120564
rect 436858 120328 436920 120564
rect 436560 120272 436920 120328
rect 438272 120564 438620 120620
rect 438272 120328 438328 120564
rect 438564 120328 438620 120564
rect 438272 120272 438620 120328
rect -23776 109694 607700 109726
rect -23776 109458 -23744 109694
rect -23508 109458 -23424 109694
rect -23188 109458 607112 109694
rect 607348 109458 607432 109694
rect 607668 109458 607700 109694
rect -23776 109374 607700 109458
rect -23776 109138 -23744 109374
rect -23508 109138 -23424 109374
rect -23188 109138 607112 109374
rect 607348 109138 607432 109374
rect 607668 109138 607700 109374
rect -23776 109106 607700 109138
rect -23776 105974 607700 106006
rect -23776 105738 -20634 105974
rect -20398 105738 -20314 105974
rect -20078 105738 604002 105974
rect 604238 105738 604322 105974
rect 604558 105738 607700 105974
rect -23776 105654 607700 105738
rect -23776 105418 -20634 105654
rect -20398 105418 -20314 105654
rect -20078 105418 604002 105654
rect 604238 105418 604322 105654
rect 604558 105418 607700 105654
rect -23776 105386 607700 105418
rect -23776 102254 607700 102286
rect -23776 102018 -17524 102254
rect -17288 102018 -17204 102254
rect -16968 102018 580626 102254
rect 580862 102018 580946 102254
rect 581182 102018 600892 102254
rect 601128 102018 601212 102254
rect 601448 102018 607700 102254
rect -23776 101934 607700 102018
rect -23776 101698 -17524 101934
rect -17288 101698 -17204 101934
rect -16968 101698 580626 101934
rect 580862 101698 580946 101934
rect 581182 101698 600892 101934
rect 601128 101698 601212 101934
rect 601448 101698 607700 101934
rect -23776 101666 607700 101698
rect -23776 98534 607700 98566
rect -23776 98298 -14414 98534
rect -14178 98298 -14094 98534
rect -13858 98298 597782 98534
rect 598018 98298 598102 98534
rect 598338 98298 607700 98534
rect -23776 98214 607700 98298
rect -23776 97978 -14414 98214
rect -14178 97978 -14094 98214
rect -13858 97978 597782 98214
rect 598018 97978 598102 98214
rect 598338 97978 607700 98214
rect -23776 97946 607700 97978
rect -23776 94814 607700 94846
rect -23776 94578 -11304 94814
rect -11068 94578 -10984 94814
rect -10748 94578 594672 94814
rect 594908 94578 594992 94814
rect 595228 94578 607700 94814
rect -23776 94494 607700 94578
rect -23776 94258 -11304 94494
rect -11068 94258 -10984 94494
rect -10748 94258 594672 94494
rect 594908 94258 594992 94494
rect 595228 94258 607700 94494
rect -23776 94226 607700 94258
rect -23776 91094 607700 91126
rect -23776 90858 -8194 91094
rect -7958 90858 -7874 91094
rect -7638 90858 591562 91094
rect 591798 90858 591882 91094
rect 592118 90858 607700 91094
rect -23776 90774 607700 90858
rect -23776 90538 -8194 90774
rect -7958 90538 -7874 90774
rect -7638 90538 591562 90774
rect 591798 90538 591882 90774
rect 592118 90538 607700 90774
rect -23776 90506 607700 90538
rect -23776 87374 607700 87406
rect -23776 87138 -5084 87374
rect -4848 87138 -4764 87374
rect -4528 87138 7876 87374
rect 8112 87138 8196 87374
rect 8432 87138 38032 87374
rect 38268 87138 38352 87374
rect 38588 87138 60622 87374
rect 60858 87138 159098 87374
rect 159334 87138 182032 87374
rect 182268 87138 182352 87374
rect 182588 87138 185622 87374
rect 185858 87138 284098 87374
rect 284334 87138 290032 87374
rect 290268 87138 290352 87374
rect 290588 87138 310622 87374
rect 310858 87138 409098 87374
rect 409334 87138 434032 87374
rect 434268 87138 434352 87374
rect 434588 87138 436622 87374
rect 436858 87138 535098 87374
rect 535334 87138 542032 87374
rect 542268 87138 542352 87374
rect 542588 87138 571532 87374
rect 571768 87138 571852 87374
rect 572088 87138 588452 87374
rect 588688 87138 588772 87374
rect 589008 87138 607700 87374
rect -23776 87054 607700 87138
rect -23776 86818 -5084 87054
rect -4848 86818 -4764 87054
rect -4528 86818 7876 87054
rect 8112 86818 8196 87054
rect 8432 86818 38032 87054
rect 38268 86818 38352 87054
rect 38588 86818 60622 87054
rect 60858 86818 159098 87054
rect 159334 86818 182032 87054
rect 182268 86818 182352 87054
rect 182588 86818 185622 87054
rect 185858 86818 284098 87054
rect 284334 86818 290032 87054
rect 290268 86818 290352 87054
rect 290588 86818 310622 87054
rect 310858 86818 409098 87054
rect 409334 86818 434032 87054
rect 434268 86818 434352 87054
rect 434588 86818 436622 87054
rect 436858 86818 535098 87054
rect 535334 86818 542032 87054
rect 542268 86818 542352 87054
rect 542588 86818 571532 87054
rect 571768 86818 571852 87054
rect 572088 86818 588452 87054
rect 588688 86818 588772 87054
rect 589008 86818 607700 87054
rect -23776 86786 607700 86818
rect -23776 83654 607700 83686
rect -23776 83418 -1974 83654
rect -1738 83418 -1654 83654
rect -1418 83418 9116 83654
rect 9352 83418 9436 83654
rect 9672 83418 56652 83654
rect 56888 83418 56972 83654
rect 57208 83418 61342 83654
rect 61578 83418 158378 83654
rect 158614 83418 164652 83654
rect 164888 83418 164972 83654
rect 165208 83418 186342 83654
rect 186578 83418 283378 83654
rect 283614 83418 308652 83654
rect 308888 83418 308972 83654
rect 309208 83418 311342 83654
rect 311578 83418 408378 83654
rect 408614 83418 416652 83654
rect 416888 83418 416972 83654
rect 417208 83418 437342 83654
rect 437578 83418 534378 83654
rect 534614 83418 560652 83654
rect 560888 83418 560972 83654
rect 561208 83418 570292 83654
rect 570528 83418 570612 83654
rect 570848 83418 585342 83654
rect 585578 83418 585662 83654
rect 585898 83418 607700 83654
rect -23776 83334 607700 83418
rect -23776 83098 -1974 83334
rect -1738 83098 -1654 83334
rect -1418 83098 9116 83334
rect 9352 83098 9436 83334
rect 9672 83098 56652 83334
rect 56888 83098 56972 83334
rect 57208 83098 61342 83334
rect 61578 83098 158378 83334
rect 158614 83098 164652 83334
rect 164888 83098 164972 83334
rect 165208 83098 186342 83334
rect 186578 83098 283378 83334
rect 283614 83098 308652 83334
rect 308888 83098 308972 83334
rect 309208 83098 311342 83334
rect 311578 83098 408378 83334
rect 408614 83098 416652 83334
rect 416888 83098 416972 83334
rect 417208 83098 437342 83334
rect 437578 83098 534378 83334
rect 534614 83098 560652 83334
rect 560888 83098 560972 83334
rect 561208 83098 570292 83334
rect 570528 83098 570612 83334
rect 570848 83098 585342 83334
rect 585578 83098 585662 83334
rect 585898 83098 607700 83334
rect -23776 83066 607700 83098
rect -23776 69694 607700 69726
rect -23776 69458 -23744 69694
rect -23508 69458 -23424 69694
rect -23188 69458 607112 69694
rect 607348 69458 607432 69694
rect 607668 69458 607700 69694
rect -23776 69374 607700 69458
rect -23776 69138 -23744 69374
rect -23508 69138 -23424 69374
rect -23188 69138 607112 69374
rect 607348 69138 607432 69374
rect 607668 69138 607700 69374
rect -23776 69106 607700 69138
rect -23776 65974 607700 66006
rect -23776 65738 -20634 65974
rect -20398 65738 -20314 65974
rect -20078 65738 604002 65974
rect 604238 65738 604322 65974
rect 604558 65738 607700 65974
rect -23776 65654 607700 65738
rect -23776 65418 -20634 65654
rect -20398 65418 -20314 65654
rect -20078 65418 604002 65654
rect 604238 65418 604322 65654
rect 604558 65418 607700 65654
rect -23776 65386 607700 65418
rect -23776 62254 607700 62286
rect -23776 62018 -17524 62254
rect -17288 62018 -17204 62254
rect -16968 62018 580626 62254
rect 580862 62018 580946 62254
rect 581182 62018 600892 62254
rect 601128 62018 601212 62254
rect 601448 62018 607700 62254
rect -23776 61934 607700 62018
rect -23776 61698 -17524 61934
rect -17288 61698 -17204 61934
rect -16968 61698 580626 61934
rect 580862 61698 580946 61934
rect 581182 61698 600892 61934
rect 601128 61698 601212 61934
rect 601448 61698 607700 61934
rect -23776 61666 607700 61698
rect -23776 58534 607700 58566
rect -23776 58298 -14414 58534
rect -14178 58298 -14094 58534
rect -13858 58298 597782 58534
rect 598018 58298 598102 58534
rect 598338 58298 607700 58534
rect -23776 58214 607700 58298
rect -23776 57978 -14414 58214
rect -14178 57978 -14094 58214
rect -13858 57978 597782 58214
rect 598018 57978 598102 58214
rect 598338 57978 607700 58214
rect -23776 57946 607700 57978
rect -23776 54814 607700 54846
rect -23776 54578 -11304 54814
rect -11068 54578 -10984 54814
rect -10748 54578 594672 54814
rect 594908 54578 594992 54814
rect 595228 54578 607700 54814
rect -23776 54494 607700 54578
rect -23776 54258 -11304 54494
rect -11068 54258 -10984 54494
rect -10748 54258 594672 54494
rect 594908 54258 594992 54494
rect 595228 54258 607700 54494
rect -23776 54226 607700 54258
rect -23776 51094 607700 51126
rect -23776 50858 -8194 51094
rect -7958 50858 -7874 51094
rect -7638 50858 591562 51094
rect 591798 50858 591882 51094
rect 592118 50858 607700 51094
rect -23776 50774 607700 50858
rect -23776 50538 -8194 50774
rect -7958 50538 -7874 50774
rect -7638 50538 591562 50774
rect 591798 50538 591882 50774
rect 592118 50538 607700 50774
rect -23776 50506 607700 50538
rect -23776 47374 607700 47406
rect -23776 47138 -5084 47374
rect -4848 47138 -4764 47374
rect -4528 47138 7876 47374
rect 8112 47138 8196 47374
rect 8432 47138 38032 47374
rect 38268 47138 38352 47374
rect 38588 47138 60622 47374
rect 60858 47138 159098 47374
rect 159334 47138 182032 47374
rect 182268 47138 182352 47374
rect 182588 47138 185622 47374
rect 185858 47138 284098 47374
rect 284334 47138 290032 47374
rect 290268 47138 290352 47374
rect 290588 47138 310622 47374
rect 310858 47138 409098 47374
rect 409334 47138 434032 47374
rect 434268 47138 434352 47374
rect 434588 47138 436622 47374
rect 436858 47138 535098 47374
rect 535334 47138 542032 47374
rect 542268 47138 542352 47374
rect 542588 47138 571532 47374
rect 571768 47138 571852 47374
rect 572088 47138 588452 47374
rect 588688 47138 588772 47374
rect 589008 47138 607700 47374
rect -23776 47054 607700 47138
rect -23776 46818 -5084 47054
rect -4848 46818 -4764 47054
rect -4528 46818 7876 47054
rect 8112 46818 8196 47054
rect 8432 46818 38032 47054
rect 38268 46818 38352 47054
rect 38588 46818 60622 47054
rect 60858 46818 159098 47054
rect 159334 46818 182032 47054
rect 182268 46818 182352 47054
rect 182588 46818 185622 47054
rect 185858 46818 284098 47054
rect 284334 46818 290032 47054
rect 290268 46818 290352 47054
rect 290588 46818 310622 47054
rect 310858 46818 409098 47054
rect 409334 46818 434032 47054
rect 434268 46818 434352 47054
rect 434588 46818 436622 47054
rect 436858 46818 535098 47054
rect 535334 46818 542032 47054
rect 542268 46818 542352 47054
rect 542588 46818 571532 47054
rect 571768 46818 571852 47054
rect 572088 46818 588452 47054
rect 588688 46818 588772 47054
rect 589008 46818 607700 47054
rect -23776 46786 607700 46818
rect -23776 43654 607700 43686
rect -23776 43418 -1974 43654
rect -1738 43418 -1654 43654
rect -1418 43418 9116 43654
rect 9352 43418 9436 43654
rect 9672 43418 56652 43654
rect 56888 43418 56972 43654
rect 57208 43418 61342 43654
rect 61578 43418 158378 43654
rect 158614 43418 164652 43654
rect 164888 43418 164972 43654
rect 165208 43418 186342 43654
rect 186578 43418 283378 43654
rect 283614 43418 308652 43654
rect 308888 43418 308972 43654
rect 309208 43418 311342 43654
rect 311578 43418 408378 43654
rect 408614 43418 416652 43654
rect 416888 43418 416972 43654
rect 417208 43418 437342 43654
rect 437578 43418 534378 43654
rect 534614 43418 560652 43654
rect 560888 43418 560972 43654
rect 561208 43418 570292 43654
rect 570528 43418 570612 43654
rect 570848 43418 585342 43654
rect 585578 43418 585662 43654
rect 585898 43418 607700 43654
rect -23776 43334 607700 43418
rect -23776 43098 -1974 43334
rect -1738 43098 -1654 43334
rect -1418 43098 9116 43334
rect 9352 43098 9436 43334
rect 9672 43098 56652 43334
rect 56888 43098 56972 43334
rect 57208 43098 61342 43334
rect 61578 43098 158378 43334
rect 158614 43098 164652 43334
rect 164888 43098 164972 43334
rect 165208 43098 186342 43334
rect 186578 43098 283378 43334
rect 283614 43098 308652 43334
rect 308888 43098 308972 43334
rect 309208 43098 311342 43334
rect 311578 43098 408378 43334
rect 408614 43098 416652 43334
rect 416888 43098 416972 43334
rect 417208 43098 437342 43334
rect 437578 43098 534378 43334
rect 534614 43098 560652 43334
rect 560888 43098 560972 43334
rect 561208 43098 570292 43334
rect 570528 43098 570612 43334
rect 570848 43098 585342 43334
rect 585578 43098 585662 43334
rect 585898 43098 607700 43334
rect -23776 43066 607700 43098
rect -23776 29694 607700 29726
rect -23776 29458 -23744 29694
rect -23508 29458 -23424 29694
rect -23188 29458 607112 29694
rect 607348 29458 607432 29694
rect 607668 29458 607700 29694
rect -23776 29374 607700 29458
rect -23776 29138 -23744 29374
rect -23508 29138 -23424 29374
rect -23188 29138 607112 29374
rect 607348 29138 607432 29374
rect 607668 29138 607700 29374
rect -23776 29106 607700 29138
rect -23776 25974 607700 26006
rect -23776 25738 -20634 25974
rect -20398 25738 -20314 25974
rect -20078 25738 604002 25974
rect 604238 25738 604322 25974
rect 604558 25738 607700 25974
rect -23776 25654 607700 25738
rect -23776 25418 -20634 25654
rect -20398 25418 -20314 25654
rect -20078 25418 604002 25654
rect 604238 25418 604322 25654
rect 604558 25418 607700 25654
rect -23776 25386 607700 25418
rect -23776 22254 607700 22286
rect -23776 22018 -17524 22254
rect -17288 22018 -17204 22254
rect -16968 22018 580626 22254
rect 580862 22018 580946 22254
rect 581182 22018 600892 22254
rect 601128 22018 601212 22254
rect 601448 22018 607700 22254
rect -23776 21934 607700 22018
rect -23776 21698 -17524 21934
rect -17288 21698 -17204 21934
rect -16968 21698 580626 21934
rect 580862 21698 580946 21934
rect 581182 21698 600892 21934
rect 601128 21698 601212 21934
rect 601448 21698 607700 21934
rect -23776 21666 607700 21698
rect 61280 21244 61640 21300
rect 61280 21008 61342 21244
rect 61578 21008 61640 21244
rect 61280 20952 61640 21008
rect 62952 21244 63300 21300
rect 62952 21008 63008 21244
rect 63244 21008 63300 21244
rect 62952 20952 63300 21008
rect 187952 21244 188300 21300
rect 187952 21008 188008 21244
rect 188244 21008 188300 21244
rect 187952 20952 188300 21008
rect 311280 21244 311640 21300
rect 311280 21008 311342 21244
rect 311578 21008 311640 21244
rect 311280 20952 311640 21008
rect 312952 21244 313300 21300
rect 312952 21008 313008 21244
rect 313244 21008 313300 21244
rect 312952 20952 313300 21008
rect 438952 21244 439300 21300
rect 438952 21008 439008 21244
rect 439244 21008 439300 21244
rect 438952 20952 439300 21008
rect 62272 20564 62620 20620
rect 62272 20328 62328 20564
rect 62564 20328 62620 20564
rect 62272 20272 62620 20328
rect 185560 20564 185920 20620
rect 185560 20328 185622 20564
rect 185858 20328 185920 20564
rect 185560 20272 185920 20328
rect 187272 20564 187620 20620
rect 187272 20328 187328 20564
rect 187564 20328 187620 20564
rect 187272 20272 187620 20328
rect 312272 20564 312620 20620
rect 312272 20328 312328 20564
rect 312564 20328 312620 20564
rect 312272 20272 312620 20328
rect 436560 20564 436920 20620
rect 436560 20328 436622 20564
rect 436858 20328 436920 20564
rect 436560 20272 436920 20328
rect 438272 20564 438620 20620
rect 438272 20328 438328 20564
rect 438564 20328 438620 20564
rect 438272 20272 438620 20328
rect 62272 19834 62620 19858
rect 62272 19598 62328 19834
rect 62564 19598 62620 19834
rect 312272 19834 312620 19858
rect 62272 19574 62620 19598
rect 187952 19578 188300 19640
rect 187952 19342 188008 19578
rect 188244 19342 188300 19578
rect 312272 19598 312328 19834
rect 312564 19598 312620 19834
rect 312272 19574 312620 19598
rect 438952 19578 439300 19640
rect 187952 19280 188300 19342
rect 438952 19342 439008 19578
rect 439244 19342 439300 19578
rect 438952 19280 439300 19342
rect -23776 18534 607700 18566
rect -23776 18298 -14414 18534
rect -14178 18298 -14094 18534
rect -13858 18298 597782 18534
rect 598018 18298 598102 18534
rect 598338 18298 607700 18534
rect -23776 18214 607700 18298
rect -23776 17978 -14414 18214
rect -14178 17978 -14094 18214
rect -13858 17978 597782 18214
rect 598018 17978 598102 18214
rect 598338 17978 607700 18214
rect -23776 17946 607700 17978
rect -23776 14814 607700 14846
rect -23776 14578 -11304 14814
rect -11068 14578 -10984 14814
rect -10748 14578 594672 14814
rect 594908 14578 594992 14814
rect 595228 14578 607700 14814
rect -23776 14494 607700 14578
rect -23776 14258 -11304 14494
rect -11068 14258 -10984 14494
rect -10748 14258 594672 14494
rect 594908 14258 594992 14494
rect 595228 14258 607700 14494
rect -23776 14226 607700 14258
rect -23776 11094 607700 11126
rect -23776 10858 -8194 11094
rect -7958 10858 -7874 11094
rect -7638 10858 591562 11094
rect 591798 10858 591882 11094
rect 592118 10858 607700 11094
rect -23776 10774 607700 10858
rect -23776 10538 -8194 10774
rect -7958 10538 -7874 10774
rect -7638 10538 591562 10774
rect 591798 10538 591882 10774
rect 592118 10538 607700 10774
rect -23776 10506 607700 10538
rect 9092 9680 9696 9712
rect 9092 9444 9116 9680
rect 9352 9444 9436 9680
rect 9672 9444 9696 9680
rect 9092 9360 9696 9444
rect 9092 9124 9116 9360
rect 9352 9124 9436 9360
rect 9672 9124 9696 9360
rect 9092 9092 9696 9124
rect 56628 9680 57232 9712
rect 56628 9444 56652 9680
rect 56888 9444 56972 9680
rect 57208 9444 57232 9680
rect 56628 9360 57232 9444
rect 56628 9124 56652 9360
rect 56888 9124 56972 9360
rect 57208 9124 57232 9360
rect 56628 9092 57232 9124
rect 92628 9680 93232 9712
rect 92628 9444 92652 9680
rect 92888 9444 92972 9680
rect 93208 9444 93232 9680
rect 92628 9360 93232 9444
rect 92628 9124 92652 9360
rect 92888 9124 92972 9360
rect 93208 9124 93232 9360
rect 92628 9092 93232 9124
rect 128628 9680 129232 9712
rect 128628 9444 128652 9680
rect 128888 9444 128972 9680
rect 129208 9444 129232 9680
rect 128628 9360 129232 9444
rect 128628 9124 128652 9360
rect 128888 9124 128972 9360
rect 129208 9124 129232 9360
rect 128628 9092 129232 9124
rect 164628 9680 165232 9712
rect 164628 9444 164652 9680
rect 164888 9444 164972 9680
rect 165208 9444 165232 9680
rect 164628 9360 165232 9444
rect 164628 9124 164652 9360
rect 164888 9124 164972 9360
rect 165208 9124 165232 9360
rect 164628 9092 165232 9124
rect 200628 9680 201232 9712
rect 200628 9444 200652 9680
rect 200888 9444 200972 9680
rect 201208 9444 201232 9680
rect 200628 9360 201232 9444
rect 200628 9124 200652 9360
rect 200888 9124 200972 9360
rect 201208 9124 201232 9360
rect 200628 9092 201232 9124
rect 236628 9680 237232 9712
rect 236628 9444 236652 9680
rect 236888 9444 236972 9680
rect 237208 9444 237232 9680
rect 236628 9360 237232 9444
rect 236628 9124 236652 9360
rect 236888 9124 236972 9360
rect 237208 9124 237232 9360
rect 236628 9092 237232 9124
rect 272628 9680 273232 9712
rect 272628 9444 272652 9680
rect 272888 9444 272972 9680
rect 273208 9444 273232 9680
rect 272628 9360 273232 9444
rect 272628 9124 272652 9360
rect 272888 9124 272972 9360
rect 273208 9124 273232 9360
rect 272628 9092 273232 9124
rect 308628 9680 309232 9712
rect 308628 9444 308652 9680
rect 308888 9444 308972 9680
rect 309208 9444 309232 9680
rect 308628 9360 309232 9444
rect 308628 9124 308652 9360
rect 308888 9124 308972 9360
rect 309208 9124 309232 9360
rect 308628 9092 309232 9124
rect 344628 9680 345232 9712
rect 344628 9444 344652 9680
rect 344888 9444 344972 9680
rect 345208 9444 345232 9680
rect 344628 9360 345232 9444
rect 344628 9124 344652 9360
rect 344888 9124 344972 9360
rect 345208 9124 345232 9360
rect 344628 9092 345232 9124
rect 380628 9680 381232 9712
rect 380628 9444 380652 9680
rect 380888 9444 380972 9680
rect 381208 9444 381232 9680
rect 380628 9360 381232 9444
rect 380628 9124 380652 9360
rect 380888 9124 380972 9360
rect 381208 9124 381232 9360
rect 380628 9092 381232 9124
rect 416628 9680 417232 9712
rect 416628 9444 416652 9680
rect 416888 9444 416972 9680
rect 417208 9444 417232 9680
rect 416628 9360 417232 9444
rect 416628 9124 416652 9360
rect 416888 9124 416972 9360
rect 417208 9124 417232 9360
rect 416628 9092 417232 9124
rect 452628 9680 453232 9712
rect 452628 9444 452652 9680
rect 452888 9444 452972 9680
rect 453208 9444 453232 9680
rect 452628 9360 453232 9444
rect 452628 9124 452652 9360
rect 452888 9124 452972 9360
rect 453208 9124 453232 9360
rect 452628 9092 453232 9124
rect 488628 9680 489232 9712
rect 488628 9444 488652 9680
rect 488888 9444 488972 9680
rect 489208 9444 489232 9680
rect 488628 9360 489232 9444
rect 488628 9124 488652 9360
rect 488888 9124 488972 9360
rect 489208 9124 489232 9360
rect 488628 9092 489232 9124
rect 524628 9680 525232 9712
rect 524628 9444 524652 9680
rect 524888 9444 524972 9680
rect 525208 9444 525232 9680
rect 524628 9360 525232 9444
rect 524628 9124 524652 9360
rect 524888 9124 524972 9360
rect 525208 9124 525232 9360
rect 524628 9092 525232 9124
rect 560628 9680 561232 9712
rect 560628 9444 560652 9680
rect 560888 9444 560972 9680
rect 561208 9444 561232 9680
rect 560628 9360 561232 9444
rect 560628 9124 560652 9360
rect 560888 9124 560972 9360
rect 561208 9124 561232 9360
rect 560628 9092 561232 9124
rect 570268 9680 570872 9712
rect 570268 9444 570292 9680
rect 570528 9444 570612 9680
rect 570848 9444 570872 9680
rect 570268 9360 570872 9444
rect 570268 9124 570292 9360
rect 570528 9124 570612 9360
rect 570848 9124 570872 9360
rect 570268 9092 570872 9124
rect 7852 8440 8456 8472
rect 7852 8204 7876 8440
rect 8112 8204 8196 8440
rect 8432 8204 8456 8440
rect 7852 8120 8456 8204
rect 7852 7884 7876 8120
rect 8112 7884 8196 8120
rect 8432 7884 8456 8120
rect 7852 7852 8456 7884
rect 38008 8440 38612 8472
rect 38008 8204 38032 8440
rect 38268 8204 38352 8440
rect 38588 8204 38612 8440
rect 38008 8120 38612 8204
rect 38008 7884 38032 8120
rect 38268 7884 38352 8120
rect 38588 7884 38612 8120
rect 38008 7852 38612 7884
rect 74008 8440 74612 8472
rect 74008 8204 74032 8440
rect 74268 8204 74352 8440
rect 74588 8204 74612 8440
rect 74008 8120 74612 8204
rect 74008 7884 74032 8120
rect 74268 7884 74352 8120
rect 74588 7884 74612 8120
rect 74008 7852 74612 7884
rect 110008 8440 110612 8472
rect 110008 8204 110032 8440
rect 110268 8204 110352 8440
rect 110588 8204 110612 8440
rect 110008 8120 110612 8204
rect 110008 7884 110032 8120
rect 110268 7884 110352 8120
rect 110588 7884 110612 8120
rect 110008 7852 110612 7884
rect 146008 8440 146612 8472
rect 146008 8204 146032 8440
rect 146268 8204 146352 8440
rect 146588 8204 146612 8440
rect 146008 8120 146612 8204
rect 146008 7884 146032 8120
rect 146268 7884 146352 8120
rect 146588 7884 146612 8120
rect 146008 7852 146612 7884
rect 182008 8440 182612 8472
rect 182008 8204 182032 8440
rect 182268 8204 182352 8440
rect 182588 8204 182612 8440
rect 182008 8120 182612 8204
rect 182008 7884 182032 8120
rect 182268 7884 182352 8120
rect 182588 7884 182612 8120
rect 182008 7852 182612 7884
rect 218008 8440 218612 8472
rect 218008 8204 218032 8440
rect 218268 8204 218352 8440
rect 218588 8204 218612 8440
rect 218008 8120 218612 8204
rect 218008 7884 218032 8120
rect 218268 7884 218352 8120
rect 218588 7884 218612 8120
rect 218008 7852 218612 7884
rect 254008 8440 254612 8472
rect 254008 8204 254032 8440
rect 254268 8204 254352 8440
rect 254588 8204 254612 8440
rect 254008 8120 254612 8204
rect 254008 7884 254032 8120
rect 254268 7884 254352 8120
rect 254588 7884 254612 8120
rect 254008 7852 254612 7884
rect 290008 8440 290612 8472
rect 290008 8204 290032 8440
rect 290268 8204 290352 8440
rect 290588 8204 290612 8440
rect 290008 8120 290612 8204
rect 290008 7884 290032 8120
rect 290268 7884 290352 8120
rect 290588 7884 290612 8120
rect 290008 7852 290612 7884
rect 326008 8440 326612 8472
rect 326008 8204 326032 8440
rect 326268 8204 326352 8440
rect 326588 8204 326612 8440
rect 326008 8120 326612 8204
rect 326008 7884 326032 8120
rect 326268 7884 326352 8120
rect 326588 7884 326612 8120
rect 326008 7852 326612 7884
rect 362008 8440 362612 8472
rect 362008 8204 362032 8440
rect 362268 8204 362352 8440
rect 362588 8204 362612 8440
rect 362008 8120 362612 8204
rect 362008 7884 362032 8120
rect 362268 7884 362352 8120
rect 362588 7884 362612 8120
rect 362008 7852 362612 7884
rect 398008 8440 398612 8472
rect 398008 8204 398032 8440
rect 398268 8204 398352 8440
rect 398588 8204 398612 8440
rect 398008 8120 398612 8204
rect 398008 7884 398032 8120
rect 398268 7884 398352 8120
rect 398588 7884 398612 8120
rect 398008 7852 398612 7884
rect 434008 8440 434612 8472
rect 434008 8204 434032 8440
rect 434268 8204 434352 8440
rect 434588 8204 434612 8440
rect 434008 8120 434612 8204
rect 434008 7884 434032 8120
rect 434268 7884 434352 8120
rect 434588 7884 434612 8120
rect 434008 7852 434612 7884
rect 470008 8440 470612 8472
rect 470008 8204 470032 8440
rect 470268 8204 470352 8440
rect 470588 8204 470612 8440
rect 470008 8120 470612 8204
rect 470008 7884 470032 8120
rect 470268 7884 470352 8120
rect 470588 7884 470612 8120
rect 470008 7852 470612 7884
rect 506008 8440 506612 8472
rect 506008 8204 506032 8440
rect 506268 8204 506352 8440
rect 506588 8204 506612 8440
rect 506008 8120 506612 8204
rect 506008 7884 506032 8120
rect 506268 7884 506352 8120
rect 506588 7884 506612 8120
rect 506008 7852 506612 7884
rect 542008 8440 542612 8472
rect 542008 8204 542032 8440
rect 542268 8204 542352 8440
rect 542588 8204 542612 8440
rect 542008 8120 542612 8204
rect 542008 7884 542032 8120
rect 542268 7884 542352 8120
rect 542588 7884 542612 8120
rect 542008 7852 542612 7884
rect 571508 8440 572112 8472
rect 571508 8204 571532 8440
rect 571768 8204 571852 8440
rect 572088 8204 572112 8440
rect 571508 8120 572112 8204
rect 571508 7884 571532 8120
rect 571768 7884 571852 8120
rect 572088 7884 572112 8120
rect 571508 7852 572112 7884
rect -23776 7374 607700 7406
rect -23776 7138 -5084 7374
rect -4848 7138 -4764 7374
rect -4528 7138 7876 7374
rect 8112 7138 8196 7374
rect 8432 7138 571532 7374
rect 571768 7138 571852 7374
rect 572088 7138 588452 7374
rect 588688 7138 588772 7374
rect 589008 7138 607700 7374
rect -23776 7054 607700 7138
rect -23776 6818 -5084 7054
rect -4848 6818 -4764 7054
rect -4528 6818 7876 7054
rect 8112 6818 8196 7054
rect 8432 6818 571532 7054
rect 571768 6818 571852 7054
rect 572088 6818 588452 7054
rect 588688 6818 588772 7054
rect 589008 6818 607700 7054
rect -23776 6786 607700 6818
rect -23776 3654 607700 3686
rect -23776 3418 -1974 3654
rect -1738 3418 -1654 3654
rect -1418 3418 585342 3654
rect 585578 3418 585662 3654
rect 585898 3418 607700 3654
rect -23776 3334 607700 3418
rect -23776 3098 -1974 3334
rect -1738 3098 -1654 3334
rect -1418 3098 585342 3334
rect 585578 3098 585662 3334
rect 585898 3098 607700 3334
rect -23776 3066 607700 3098
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -5116 -3456 589040 -3424
rect -5116 -3692 -5084 -3456
rect -4848 -3692 -4764 -3456
rect -4528 -3692 588452 -3456
rect 588688 -3692 588772 -3456
rect 589008 -3692 589040 -3456
rect -5116 -3776 589040 -3692
rect -5116 -4012 -5084 -3776
rect -4848 -4012 -4764 -3776
rect -4528 -4012 588452 -3776
rect 588688 -4012 588772 -3776
rect 589008 -4012 589040 -3776
rect -5116 -4044 589040 -4012
rect -8226 -6566 592150 -6534
rect -8226 -6802 -8194 -6566
rect -7958 -6802 -7874 -6566
rect -7638 -6802 591562 -6566
rect 591798 -6802 591882 -6566
rect 592118 -6802 592150 -6566
rect -8226 -6886 592150 -6802
rect -8226 -7122 -8194 -6886
rect -7958 -7122 -7874 -6886
rect -7638 -7122 591562 -6886
rect 591798 -7122 591882 -6886
rect 592118 -7122 592150 -6886
rect -8226 -7154 592150 -7122
rect -11336 -9676 595260 -9644
rect -11336 -9912 -11304 -9676
rect -11068 -9912 -10984 -9676
rect -10748 -9912 594672 -9676
rect 594908 -9912 594992 -9676
rect 595228 -9912 595260 -9676
rect -11336 -9996 595260 -9912
rect -11336 -10232 -11304 -9996
rect -11068 -10232 -10984 -9996
rect -10748 -10232 594672 -9996
rect 594908 -10232 594992 -9996
rect 595228 -10232 595260 -9996
rect -11336 -10264 595260 -10232
rect -14446 -12786 598370 -12754
rect -14446 -13022 -14414 -12786
rect -14178 -13022 -14094 -12786
rect -13858 -13022 597782 -12786
rect 598018 -13022 598102 -12786
rect 598338 -13022 598370 -12786
rect -14446 -13106 598370 -13022
rect -14446 -13342 -14414 -13106
rect -14178 -13342 -14094 -13106
rect -13858 -13342 597782 -13106
rect 598018 -13342 598102 -13106
rect 598338 -13342 598370 -13106
rect -14446 -13374 598370 -13342
rect -17556 -15896 601480 -15864
rect -17556 -16132 -17524 -15896
rect -17288 -16132 -17204 -15896
rect -16968 -16132 580626 -15896
rect 580862 -16132 580946 -15896
rect 581182 -16132 600892 -15896
rect 601128 -16132 601212 -15896
rect 601448 -16132 601480 -15896
rect -17556 -16216 601480 -16132
rect -17556 -16452 -17524 -16216
rect -17288 -16452 -17204 -16216
rect -16968 -16452 580626 -16216
rect 580862 -16452 580946 -16216
rect 581182 -16452 600892 -16216
rect 601128 -16452 601212 -16216
rect 601448 -16452 601480 -16216
rect -17556 -16484 601480 -16452
rect -20666 -19006 604590 -18974
rect -20666 -19242 -20634 -19006
rect -20398 -19242 -20314 -19006
rect -20078 -19242 604002 -19006
rect 604238 -19242 604322 -19006
rect 604558 -19242 604590 -19006
rect -20666 -19326 604590 -19242
rect -20666 -19562 -20634 -19326
rect -20398 -19562 -20314 -19326
rect -20078 -19562 604002 -19326
rect 604238 -19562 604322 -19326
rect 604558 -19562 604590 -19326
rect -20666 -19594 604590 -19562
rect -23776 -22116 607700 -22084
rect -23776 -22352 -23744 -22116
rect -23508 -22352 -23424 -22116
rect -23188 -22352 607112 -22116
rect 607348 -22352 607432 -22116
rect 607668 -22352 607700 -22116
rect -23776 -22436 607700 -22352
rect -23776 -22672 -23744 -22436
rect -23508 -22672 -23424 -22436
rect -23188 -22672 607112 -22436
rect 607348 -22672 607432 -22436
rect 607668 -22672 607700 -22436
rect -23776 -22704 607700 -22672
use user_proj_example  mprj
timestamp 0
transform 1 0 4000 0 1 4000
box 0 0 571964 694008
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 3066 607700 3686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 43066 607700 43686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 83066 607700 83686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 123066 607700 123686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 163066 607700 163686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 203066 607700 203686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 243066 607700 243686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 283066 607700 283686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 323066 607700 323686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 363066 607700 363686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 403066 607700 403686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 443066 607700 443686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 483066 607700 483686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 523066 607700 523686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 563066 607700 563686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 603066 607700 603686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 643066 607700 643686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 683066 607700 683686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -8226 -7154 -7606 711090 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8226 -7154 592150 -6534 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8226 710470 592150 711090 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 591530 -7154 592150 711090 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 10506 607700 11126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 50506 607700 51126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 90506 607700 91126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 130506 607700 131126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 170506 607700 171126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 210506 607700 211126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 250506 607700 251126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 290506 607700 291126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 330506 607700 331126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 370506 607700 371126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 410506 607700 411126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 450506 607700 451126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 490506 607700 491126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 530506 607700 531126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 570506 607700 571126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 610506 607700 611126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 650506 607700 651126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 690506 607700 691126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -14446 -13374 -13826 717310 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -14446 -13374 598370 -12754 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -14446 716690 598370 717310 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 597750 -13374 598370 717310 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 17946 607700 18566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 57946 607700 58566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 97946 607700 98566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 137946 607700 138566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 177946 607700 178566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 217946 607700 218566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 257946 607700 258566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 297946 607700 298566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 337946 607700 338566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 377946 607700 378566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 417946 607700 418566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 457946 607700 458566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 497946 607700 498566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 537946 607700 538566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 577946 607700 578566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 617946 607700 618566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 657946 607700 658566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 697946 607700 698566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -20666 -19594 -20046 723530 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -20666 -19594 604590 -18974 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -20666 722910 604590 723530 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 603970 -19594 604590 723530 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 25386 607700 26006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 65386 607700 66006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 105386 607700 106006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 145386 607700 146006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 185386 607700 186006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 225386 607700 226006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 265386 607700 266006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 305386 607700 306006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 345386 607700 346006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 385386 607700 386006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 425386 607700 426006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 465386 607700 466006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 505386 607700 506006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 545386 607700 546006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 585386 607700 586006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 625386 607700 626006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 665386 607700 666006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -17556 -16484 -16936 720420 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -17556 -16484 601480 -15864 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -17556 719800 601480 720420 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 600860 -16484 601480 720420 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 580594 -22704 581214 726640 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 21666 607700 22286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 61666 607700 62286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 101666 607700 102286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 141666 607700 142286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 181666 607700 182286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 221666 607700 222286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 261666 607700 262286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 301666 607700 302286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 341666 607700 342286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 381666 607700 382286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 421666 607700 422286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 461666 607700 462286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 501666 607700 502286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 541666 607700 542286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 581666 607700 582286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 621666 607700 622286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 661666 607700 662286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -23776 -22704 -23156 726640 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 -22704 607700 -22084 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 726020 607700 726640 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 607080 -22704 607700 726640 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 29106 607700 29726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 69106 607700 69726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 109106 607700 109726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 149106 607700 149726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 189106 607700 189726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 229106 607700 229726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 269106 607700 269726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 309106 607700 309726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 349106 607700 349726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 389106 607700 389726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 429106 607700 429726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 469106 607700 469726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 509106 607700 509726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 549106 607700 549726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 589106 607700 589726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 629106 607700 629726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 669106 607700 669726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -5116 -4044 -4496 707980 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -5116 -4044 589040 -3424 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -5116 707360 589040 707980 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 588420 -4044 589040 707980 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 6786 607700 7406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 46786 607700 47406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 86786 607700 87406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 126786 607700 127406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 166786 607700 167406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 206786 607700 207406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 246786 607700 247406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 286786 607700 287406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 326786 607700 327406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 366786 607700 367406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 406786 607700 407406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 446786 607700 447406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 486786 607700 487406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 526786 607700 527406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 566786 607700 567406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 606786 607700 607406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 646786 607700 647406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 686786 607700 687406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -11336 -10264 -10716 714200 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -11336 -10264 595260 -9644 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -11336 713580 595260 714200 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 594640 -10264 595260 714200 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 14226 607700 14846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 54226 607700 54846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 94226 607700 94846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 134226 607700 134846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 174226 607700 174846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 214226 607700 214846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 254226 607700 254846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 294226 607700 294846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 334226 607700 334846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 374226 607700 374846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 414226 607700 414846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 454226 607700 454846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 494226 607700 494846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 534226 607700 534846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 574226 607700 574846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 614226 607700 614846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 654226 607700 654846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 694226 607700 694846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
rlabel via4 570730 692358 570730 692358 0 vccd1
rlabel metal5 291962 690816 291962 690816 0 vccd2
rlabel metal5 291962 698256 291962 698256 0 vdda1
rlabel metal5 291962 665696 291962 665696 0 vdda2
rlabel metal5 291962 661976 291962 661976 0 vssa1
rlabel metal5 291962 669416 291962 669416 0 vssa2
rlabel via4 571970 693598 571970 693598 0 vssd1
rlabel metal5 291962 694536 291962 694536 0 vssd2
rlabel metal2 580198 284920 580198 284920 0 analog_io[0]
rlabel metal2 445186 698064 445186 698064 0 analog_io[10]
rlabel metal2 379774 698064 379774 698064 0 analog_io[11]
rlabel metal2 314454 698064 314454 698064 0 analog_io[12]
rlabel metal2 249042 698064 249042 698064 0 analog_io[13]
rlabel metal2 183722 698064 183722 698064 0 analog_io[14]
rlabel metal2 118402 698064 118402 698064 0 analog_io[15]
rlabel metal2 56810 702076 56810 702076 0 analog_io[16]
rlabel metal3 3780 697948 3780 697948 0 analog_io[17]
rlabel metal3 3711 645488 3711 645488 0 analog_io[18]
rlabel metal3 3711 593150 3711 593150 0 analog_io[19]
rlabel metal2 579600 337892 579600 337892 0 analog_io[1]
rlabel metal3 3711 540812 3711 540812 0 analog_io[20]
rlabel metal3 3711 488474 3711 488474 0 analog_io[21]
rlabel metal3 3734 436014 3734 436014 0 analog_io[22]
rlabel metal3 3734 383676 3734 383676 0 analog_io[23]
rlabel metal3 3734 331338 3734 331338 0 analog_io[24]
rlabel metal3 3734 279000 3734 279000 0 analog_io[25]
rlabel metal3 3734 226662 3734 226662 0 analog_io[26]
rlabel metal3 3734 174202 3734 174202 0 analog_io[27]
rlabel metal3 3734 121864 3734 121864 0 analog_io[28]
rlabel metal3 583556 391408 583556 391408 0 analog_io[2]
rlabel metal3 580183 444788 580183 444788 0 analog_io[3]
rlabel metal3 576165 497868 576165 497868 0 analog_io[4]
rlabel metal3 576165 551182 576165 551182 0 analog_io[5]
rlabel metal3 579692 604316 579692 604316 0 analog_io[6]
rlabel metal3 583556 657696 583556 657696 0 analog_io[7]
rlabel metal2 575918 698064 575918 698064 0 analog_io[8]
rlabel metal2 510506 698064 510506 698064 0 analog_io[9]
rlabel metal2 576886 4845 576886 4845 0 io_in[0]
rlabel metal3 580183 458116 580183 458116 0 io_in[10]
rlabel metal3 576165 511166 576165 511166 0 io_in[11]
rlabel metal3 579692 564400 579692 564400 0 io_in[12]
rlabel metal3 583556 617780 583556 617780 0 io_in[13]
rlabel metal3 583556 671092 583556 671092 0 io_in[14]
rlabel metal2 559542 698064 559542 698064 0 io_in[15]
rlabel metal2 494222 698064 494222 698064 0 io_in[16]
rlabel metal2 428810 698064 428810 698064 0 io_in[17]
rlabel metal2 365010 701974 365010 701974 0 io_in[18]
rlabel metal2 298078 698064 298078 698064 0 io_in[19]
rlabel metal2 578358 44625 578358 44625 0 io_in[1]
rlabel metal2 232758 698064 232758 698064 0 io_in[20]
rlabel metal2 167346 698064 167346 698064 0 io_in[21]
rlabel metal2 102026 698064 102026 698064 0 io_in[22]
rlabel metal2 36706 698064 36706 698064 0 io_in[23]
rlabel metal3 3711 684772 3711 684772 0 io_in[24]
rlabel metal3 3711 632434 3711 632434 0 io_in[25]
rlabel metal3 3711 580096 3711 580096 0 io_in[26]
rlabel metal3 3711 527758 3711 527758 0 io_in[27]
rlabel metal3 3711 475298 3711 475298 0 io_in[28]
rlabel metal3 3734 422960 3734 422960 0 io_in[29]
rlabel metal2 579600 84252 579600 84252 0 io_in[2]
rlabel metal3 3734 370622 3734 370622 0 io_in[30]
rlabel metal3 3734 318284 3734 318284 0 io_in[31]
rlabel metal3 3734 265946 3734 265946 0 io_in[32]
rlabel metal3 3734 213486 3734 213486 0 io_in[33]
rlabel metal3 3711 161148 3711 161148 0 io_in[34]
rlabel metal3 3711 108810 3711 108810 0 io_in[35]
rlabel metal3 3734 69526 3734 69526 0 io_in[36]
rlabel metal3 3711 30242 3711 30242 0 io_in[37]
rlabel metal2 579600 124372 579600 124372 0 io_in[3]
rlabel metal2 579600 164356 579600 164356 0 io_in[4]
rlabel metal2 579600 204340 579600 204340 0 io_in[5]
rlabel metal2 580198 245004 580198 245004 0 io_in[6]
rlabel metal2 579600 297772 579600 297772 0 io_in[7]
rlabel metal2 579554 351492 579554 351492 0 io_in[8]
rlabel metal3 583556 404668 583556 404668 0 io_in[9]
rlabel metal2 579600 30940 579600 30940 0 io_oeb[0]
rlabel metal3 576165 484570 576165 484570 0 io_oeb[10]
rlabel metal3 576165 537884 576165 537884 0 io_oeb[11]
rlabel metal3 580183 590988 580183 590988 0 io_oeb[12]
rlabel metal3 582230 644028 582230 644028 0 io_oeb[13]
rlabel metal2 580198 697731 580198 697731 0 io_oeb[14]
rlabel metal2 526882 698064 526882 698064 0 io_oeb[15]
rlabel metal2 461470 698064 461470 698064 0 io_oeb[16]
rlabel metal2 396150 698064 396150 698064 0 io_oeb[17]
rlabel metal2 330738 698064 330738 698064 0 io_oeb[18]
rlabel metal2 265418 698064 265418 698064 0 io_oeb[19]
rlabel metal2 579600 70924 579600 70924 0 io_oeb[1]
rlabel metal2 200098 698064 200098 698064 0 io_oeb[20]
rlabel metal2 134686 698064 134686 698064 0 io_oeb[21]
rlabel metal2 69366 698064 69366 698064 0 io_oeb[22]
rlabel metal2 4046 698081 4046 698081 0 io_oeb[23]
rlabel metal3 3711 658664 3711 658664 0 io_oeb[24]
rlabel metal3 3711 606204 3711 606204 0 io_oeb[25]
rlabel metal3 3711 553866 3711 553866 0 io_oeb[26]
rlabel metal3 3711 501528 3711 501528 0 io_oeb[27]
rlabel metal3 3711 449190 3711 449190 0 io_oeb[28]
rlabel metal3 3734 396852 3734 396852 0 io_oeb[29]
rlabel metal2 579600 110908 579600 110908 0 io_oeb[2]
rlabel metal3 1878 345372 1878 345372 0 io_oeb[30]
rlabel metal3 3734 292054 3734 292054 0 io_oeb[31]
rlabel metal3 3734 239716 3734 239716 0 io_oeb[32]
rlabel metal3 3826 187378 3826 187378 0 io_oeb[33]
rlabel metal3 3711 135040 3711 135040 0 io_oeb[34]
rlabel metal3 3711 82580 3711 82580 0 io_oeb[35]
rlabel metal3 3734 43296 3734 43296 0 io_oeb[36]
rlabel metal3 3895 4134 3895 4134 0 io_oeb[37]
rlabel metal3 582230 152660 582230 152660 0 io_oeb[3]
rlabel metal2 579600 191012 579600 191012 0 io_oeb[4]
rlabel metal2 579600 231132 579600 231132 0 io_oeb[5]
rlabel metal2 579600 271116 579600 271116 0 io_oeb[6]
rlabel metal2 580198 324836 580198 324836 0 io_oeb[7]
rlabel metal3 579508 378012 579508 378012 0 io_oeb[8]
rlabel metal3 583556 431324 583556 431324 0 io_oeb[9]
rlabel metal2 579600 17612 579600 17612 0 io_out[0]
rlabel metal3 580183 471444 580183 471444 0 io_out[10]
rlabel metal3 576165 524586 576165 524586 0 io_out[11]
rlabel metal3 580183 577660 580183 577660 0 io_out[12]
rlabel metal3 583556 631108 583556 631108 0 io_out[13]
rlabel metal2 579600 684692 579600 684692 0 io_out[14]
rlabel metal2 543166 698064 543166 698064 0 io_out[15]
rlabel metal2 477846 698064 477846 698064 0 io_out[16]
rlabel metal2 412434 698064 412434 698064 0 io_out[17]
rlabel metal2 347114 698064 347114 698064 0 io_out[18]
rlabel metal2 281794 698064 281794 698064 0 io_out[19]
rlabel metal2 579600 57596 579600 57596 0 io_out[1]
rlabel metal2 216382 698064 216382 698064 0 io_out[20]
rlabel metal2 154146 702076 154146 702076 0 io_out[21]
rlabel metal2 85742 698064 85742 698064 0 io_out[22]
rlabel metal2 20330 698064 20330 698064 0 io_out[23]
rlabel metal3 3711 671718 3711 671718 0 io_out[24]
rlabel metal3 3711 619380 3711 619380 0 io_out[25]
rlabel metal3 3711 566920 3711 566920 0 io_out[26]
rlabel metal3 3711 514582 3711 514582 0 io_out[27]
rlabel metal3 3711 462244 3711 462244 0 io_out[28]
rlabel metal3 3734 409906 3734 409906 0 io_out[29]
rlabel metal2 579600 97580 579600 97580 0 io_out[2]
rlabel metal3 3734 357568 3734 357568 0 io_out[30]
rlabel metal3 3734 305108 3734 305108 0 io_out[31]
rlabel metal3 3734 252770 3734 252770 0 io_out[32]
rlabel metal3 3734 200432 3734 200432 0 io_out[33]
rlabel metal3 3734 148094 3734 148094 0 io_out[34]
rlabel metal3 3734 95756 3734 95756 0 io_out[35]
rlabel metal3 3711 56472 3711 56472 0 io_out[36]
rlabel metal3 3711 17188 3711 17188 0 io_out[37]
rlabel metal2 579600 137564 579600 137564 0 io_out[3]
rlabel metal2 579600 177684 579600 177684 0 io_out[4]
rlabel metal2 579600 217668 579600 217668 0 io_out[5]
rlabel metal2 578910 257737 578910 257737 0 io_out[6]
rlabel metal2 579600 311100 579600 311100 0 io_out[7]
rlabel metal3 583556 364684 583556 364684 0 io_out[8]
rlabel metal3 579692 418200 579692 418200 0 io_out[9]
rlabel metal2 125902 840 125902 840 0 la_data_in[0]
rlabel metal2 480562 772 480562 772 0 la_data_in[100]
rlabel metal2 484058 1588 484058 1588 0 la_data_in[101]
rlabel metal2 487455 340 487455 340 0 la_data_in[102]
rlabel metal2 485530 2397 485530 2397 0 la_data_in[103]
rlabel metal2 489026 2499 489026 2499 0 la_data_in[104]
rlabel metal2 498226 772 498226 772 0 la_data_in[105]
rlabel metal2 501814 670 501814 670 0 la_data_in[106]
rlabel via1 505586 51 505586 51 0 la_data_in[107]
rlabel metal2 508898 670 508898 670 0 la_data_in[108]
rlabel metal2 506322 1887 506322 1887 0 la_data_in[109]
rlabel metal2 161598 2040 161598 2040 0 la_data_in[10]
rlabel metal2 515883 340 515883 340 0 la_data_in[110]
rlabel metal2 519570 772 519570 772 0 la_data_in[111]
rlabel via1 523250 51 523250 51 0 la_data_in[112]
rlabel metal2 526654 670 526654 670 0 la_data_in[113]
rlabel metal2 523802 2431 523802 2431 0 la_data_in[114]
rlabel metal2 527298 2499 527298 2499 0 la_data_in[115]
rlabel metal2 537234 738 537234 738 0 la_data_in[116]
rlabel metal2 540631 340 540631 340 0 la_data_in[117]
rlabel via1 544594 323 544594 323 0 la_data_in[118]
rlabel metal2 541190 2227 541190 2227 0 la_data_in[119]
rlabel metal2 164910 2047 164910 2047 0 la_data_in[11]
rlabel metal2 544686 2091 544686 2091 0 la_data_in[120]
rlabel metal2 554990 772 554990 772 0 la_data_in[121]
rlabel metal2 558578 840 558578 840 0 la_data_in[122]
rlabel via1 562258 85 562258 85 0 la_data_in[123]
rlabel metal2 565662 772 565662 772 0 la_data_in[124]
rlabel metal2 562074 2499 562074 2499 0 la_data_in[125]
rlabel metal2 565478 1921 565478 1921 0 la_data_in[126]
rlabel metal2 576334 772 576334 772 0 la_data_in[127]
rlabel metal2 168406 2047 168406 2047 0 la_data_in[12]
rlabel metal2 172139 340 172139 340 0 la_data_in[13]
rlabel metal2 175635 340 175635 340 0 la_data_in[14]
rlabel metal2 179078 2047 179078 2047 0 la_data_in[15]
rlabel metal2 182574 2047 182574 2047 0 la_data_in[16]
rlabel metal2 186162 2047 186162 2047 0 la_data_in[17]
rlabel metal2 189750 2047 189750 2047 0 la_data_in[18]
rlabel metal2 193246 2047 193246 2047 0 la_data_in[19]
rlabel metal2 129398 840 129398 840 0 la_data_in[1]
rlabel metal2 196834 2047 196834 2047 0 la_data_in[20]
rlabel metal2 200098 3869 200098 3869 0 la_data_in[21]
rlabel metal2 203773 340 203773 340 0 la_data_in[22]
rlabel metal2 207269 340 207269 340 0 la_data_in[23]
rlabel metal2 211002 2047 211002 2047 0 la_data_in[24]
rlabel metal2 214498 2047 214498 2047 0 la_data_in[25]
rlabel metal2 217849 340 217849 340 0 la_data_in[26]
rlabel metal2 221345 340 221345 340 0 la_data_in[27]
rlabel metal2 225170 2064 225170 2064 0 la_data_in[28]
rlabel metal2 228521 340 228521 340 0 la_data_in[29]
rlabel metal2 132986 840 132986 840 0 la_data_in[2]
rlabel metal2 232254 2064 232254 2064 0 la_data_in[30]
rlabel metal2 235842 2047 235842 2047 0 la_data_in[31]
rlabel metal2 238370 3886 238370 3886 0 la_data_in[32]
rlabel metal2 242926 2064 242926 2064 0 la_data_in[33]
rlabel metal2 246422 2064 246422 2064 0 la_data_in[34]
rlabel metal2 250010 1588 250010 1588 0 la_data_in[35]
rlabel metal2 253506 2064 253506 2064 0 la_data_in[36]
rlabel metal2 257094 2064 257094 2064 0 la_data_in[37]
rlabel metal2 260682 2098 260682 2098 0 la_data_in[38]
rlabel metal2 264178 2064 264178 2064 0 la_data_in[39]
rlabel metal2 136482 806 136482 806 0 la_data_in[3]
rlabel metal2 267766 840 267766 840 0 la_data_in[40]
rlabel metal2 271262 2064 271262 2064 0 la_data_in[41]
rlabel metal2 274850 840 274850 840 0 la_data_in[42]
rlabel metal2 276734 3886 276734 3886 0 la_data_in[43]
rlabel metal2 281934 840 281934 840 0 la_data_in[44]
rlabel metal2 285430 2064 285430 2064 0 la_data_in[45]
rlabel metal2 289018 2064 289018 2064 0 la_data_in[46]
rlabel metal2 292606 466 292606 466 0 la_data_in[47]
rlabel metal2 296102 2064 296102 2064 0 la_data_in[48]
rlabel metal2 299690 840 299690 840 0 la_data_in[49]
rlabel metal2 140070 806 140070 806 0 la_data_in[4]
rlabel metal2 303186 2064 303186 2064 0 la_data_in[50]
rlabel metal2 306774 466 306774 466 0 la_data_in[51]
rlabel metal2 310270 2064 310270 2064 0 la_data_in[52]
rlabel metal2 313858 772 313858 772 0 la_data_in[53]
rlabel metal2 315054 3281 315054 3281 0 la_data_in[54]
rlabel metal2 320942 806 320942 806 0 la_data_in[55]
rlabel metal2 324438 840 324438 840 0 la_data_in[56]
rlabel metal2 328026 840 328026 840 0 la_data_in[57]
rlabel metal2 331614 840 331614 840 0 la_data_in[58]
rlabel metal2 335110 840 335110 840 0 la_data_in[59]
rlabel metal2 143566 2047 143566 2047 0 la_data_in[5]
rlabel metal2 338698 840 338698 840 0 la_data_in[60]
rlabel metal2 342194 840 342194 840 0 la_data_in[61]
rlabel metal2 345782 534 345782 534 0 la_data_in[62]
rlabel metal2 349278 534 349278 534 0 la_data_in[63]
rlabel metal2 352866 840 352866 840 0 la_data_in[64]
rlabel metal2 353234 2533 353234 2533 0 la_data_in[65]
rlabel metal2 359950 840 359950 840 0 la_data_in[66]
rlabel metal2 363538 738 363538 738 0 la_data_in[67]
rlabel metal2 367034 806 367034 806 0 la_data_in[68]
rlabel metal2 370622 840 370622 840 0 la_data_in[69]
rlabel metal2 147391 340 147391 340 0 la_data_in[6]
rlabel metal2 370714 2533 370714 2533 0 la_data_in[70]
rlabel metal2 377706 670 377706 670 0 la_data_in[71]
rlabel metal2 381202 806 381202 806 0 la_data_in[72]
rlabel metal2 384790 772 384790 772 0 la_data_in[73]
rlabel metal2 388286 602 388286 602 0 la_data_in[74]
rlabel metal2 391874 806 391874 806 0 la_data_in[75]
rlabel metal2 391598 2295 391598 2295 0 la_data_in[76]
rlabel metal2 398958 840 398958 840 0 la_data_in[77]
rlabel metal2 402546 806 402546 806 0 la_data_in[78]
rlabel via1 406226 51 406226 51 0 la_data_in[79]
rlabel metal2 150887 340 150887 340 0 la_data_in[7]
rlabel metal2 409630 840 409630 840 0 la_data_in[80]
rlabel metal2 408986 2431 408986 2431 0 la_data_in[81]
rlabel metal2 412482 1989 412482 1989 0 la_data_in[82]
rlabel metal2 420210 840 420210 840 0 la_data_in[83]
rlabel metal2 423607 340 423607 340 0 la_data_in[84]
rlabel metal2 427294 670 427294 670 0 la_data_in[85]
rlabel metal2 430882 772 430882 772 0 la_data_in[86]
rlabel metal2 429870 2295 429870 2295 0 la_data_in[87]
rlabel metal2 437966 551 437966 551 0 la_data_in[88]
rlabel metal2 441554 738 441554 738 0 la_data_in[89]
rlabel metal2 154238 840 154238 840 0 la_data_in[8]
rlabel metal2 445050 1588 445050 1588 0 la_data_in[90]
rlabel metal2 448447 340 448447 340 0 la_data_in[91]
rlabel metal2 447258 2397 447258 2397 0 la_data_in[92]
rlabel metal2 450754 2499 450754 2499 0 la_data_in[93]
rlabel metal2 459218 738 459218 738 0 la_data_in[94]
rlabel metal2 462615 340 462615 340 0 la_data_in[95]
rlabel metal2 466302 738 466302 738 0 la_data_in[96]
rlabel metal2 469890 670 469890 670 0 la_data_in[97]
rlabel metal2 468142 2533 468142 2533 0 la_data_in[98]
rlabel metal2 476783 340 476783 340 0 la_data_in[99]
rlabel metal2 158063 340 158063 340 0 la_data_in[9]
rlabel metal2 127006 755 127006 755 0 la_data_out[0]
rlabel metal2 481567 340 481567 340 0 la_data_out[100]
rlabel metal2 485063 340 485063 340 0 la_data_out[101]
rlabel metal2 488842 636 488842 636 0 la_data_out[102]
rlabel metal2 486726 2431 486726 2431 0 la_data_out[103]
rlabel metal2 495735 340 495735 340 0 la_data_out[104]
rlabel metal2 499422 738 499422 738 0 la_data_out[105]
rlabel metal2 503010 840 503010 840 0 la_data_out[106]
rlabel metal2 506506 738 506506 738 0 la_data_out[107]
rlabel metal2 504114 2533 504114 2533 0 la_data_out[108]
rlabel metal2 507518 2091 507518 2091 0 la_data_out[109]
rlabel metal2 162518 840 162518 840 0 la_data_out[10]
rlabel metal2 517178 806 517178 806 0 la_data_out[110]
rlabel metal2 520766 704 520766 704 0 la_data_out[111]
rlabel metal2 524071 340 524071 340 0 la_data_out[112]
rlabel metal2 527850 704 527850 704 0 la_data_out[113]
rlabel metal2 524998 1921 524998 1921 0 la_data_out[114]
rlabel metal2 528494 1989 528494 1989 0 la_data_out[115]
rlabel metal2 538430 772 538430 772 0 la_data_out[116]
rlabel metal2 542117 340 542117 340 0 la_data_out[117]
rlabel metal2 545514 738 545514 738 0 la_data_out[118]
rlabel metal2 542294 2533 542294 2533 0 la_data_out[119]
rlabel metal2 166297 340 166297 340 0 la_data_out[11]
rlabel metal2 545882 2023 545882 2023 0 la_data_out[120]
rlabel metal2 556186 704 556186 704 0 la_data_out[121]
rlabel metal2 559774 738 559774 738 0 la_data_out[122]
rlabel metal2 563270 466 563270 466 0 la_data_out[123]
rlabel metal2 566858 704 566858 704 0 la_data_out[124]
rlabel metal2 563178 2193 563178 2193 0 la_data_out[125]
rlabel metal2 566674 2091 566674 2091 0 la_data_out[126]
rlabel metal2 577438 806 577438 806 0 la_data_out[127]
rlabel metal2 169793 340 169793 340 0 la_data_out[12]
rlabel metal2 173190 2047 173190 2047 0 la_data_out[13]
rlabel metal2 176686 2047 176686 2047 0 la_data_out[14]
rlabel metal2 180373 204 180373 204 0 la_data_out[15]
rlabel metal2 183869 204 183869 204 0 la_data_out[16]
rlabel metal2 187358 2047 187358 2047 0 la_data_out[17]
rlabel metal2 190854 2047 190854 2047 0 la_data_out[18]
rlabel metal2 194442 2047 194442 2047 0 la_data_out[19]
rlabel metal2 130594 840 130594 840 0 la_data_out[1]
rlabel metal2 197938 2047 197938 2047 0 la_data_out[20]
rlabel metal2 201427 340 201427 340 0 la_data_out[21]
rlabel metal2 205114 2047 205114 2047 0 la_data_out[22]
rlabel metal2 208610 2047 208610 2047 0 la_data_out[23]
rlabel metal2 211961 340 211961 340 0 la_data_out[24]
rlabel metal2 215457 340 215457 340 0 la_data_out[25]
rlabel metal2 219282 2047 219282 2047 0 la_data_out[26]
rlabel metal2 222778 2064 222778 2064 0 la_data_out[27]
rlabel metal2 226129 340 226129 340 0 la_data_out[28]
rlabel metal2 229625 340 229625 340 0 la_data_out[29]
rlabel metal2 134182 2047 134182 2047 0 la_data_out[2]
rlabel metal2 233450 2064 233450 2064 0 la_data_out[30]
rlabel metal2 236801 340 236801 340 0 la_data_out[31]
rlabel metal2 240534 2064 240534 2064 0 la_data_out[32]
rlabel metal2 244122 2047 244122 2047 0 la_data_out[33]
rlabel metal2 247618 2064 247618 2064 0 la_data_out[34]
rlabel metal2 251206 2064 251206 2064 0 la_data_out[35]
rlabel metal2 254702 1622 254702 1622 0 la_data_out[36]
rlabel metal2 256954 3920 256954 3920 0 la_data_out[37]
rlabel metal2 261786 2064 261786 2064 0 la_data_out[38]
rlabel metal2 265374 2098 265374 2098 0 la_data_out[39]
rlabel metal2 137678 840 137678 840 0 la_data_out[3]
rlabel metal2 268870 2064 268870 2064 0 la_data_out[40]
rlabel metal2 272458 2098 272458 2098 0 la_data_out[41]
rlabel metal2 276046 534 276046 534 0 la_data_out[42]
rlabel metal2 279542 2098 279542 2098 0 la_data_out[43]
rlabel metal2 283130 806 283130 806 0 la_data_out[44]
rlabel metal2 286626 2098 286626 2098 0 la_data_out[45]
rlabel metal2 290214 840 290214 840 0 la_data_out[46]
rlabel metal2 293710 2064 293710 2064 0 la_data_out[47]
rlabel metal2 295274 2533 295274 2533 0 la_data_out[48]
rlabel metal2 300794 2064 300794 2064 0 la_data_out[49]
rlabel metal2 141503 340 141503 340 0 la_data_out[4]
rlabel metal2 304382 840 304382 840 0 la_data_out[50]
rlabel metal2 307970 840 307970 840 0 la_data_out[51]
rlabel metal2 311466 1588 311466 1588 0 la_data_out[52]
rlabel metal2 315054 806 315054 806 0 la_data_out[53]
rlabel metal2 318550 2064 318550 2064 0 la_data_out[54]
rlabel metal2 322138 772 322138 772 0 la_data_out[55]
rlabel metal2 325634 2064 325634 2064 0 la_data_out[56]
rlabel metal2 329222 772 329222 772 0 la_data_out[57]
rlabel metal2 332718 806 332718 806 0 la_data_out[58]
rlabel metal2 333546 2227 333546 2227 0 la_data_out[59]
rlabel metal2 144762 840 144762 840 0 la_data_out[5]
rlabel metal2 339894 772 339894 772 0 la_data_out[60]
rlabel metal2 343390 806 343390 806 0 la_data_out[61]
rlabel metal2 346978 806 346978 806 0 la_data_out[62]
rlabel metal2 350474 602 350474 602 0 la_data_out[63]
rlabel metal2 354062 534 354062 534 0 la_data_out[64]
rlabel metal2 354430 1887 354430 1887 0 la_data_out[65]
rlabel metal2 361146 772 361146 772 0 la_data_out[66]
rlabel metal2 364642 602 364642 602 0 la_data_out[67]
rlabel metal2 368230 772 368230 772 0 la_data_out[68]
rlabel metal2 371726 602 371726 602 0 la_data_out[69]
rlabel metal2 148350 840 148350 840 0 la_data_out[6]
rlabel metal2 371818 2295 371818 2295 0 la_data_out[70]
rlabel metal2 378902 772 378902 772 0 la_data_out[71]
rlabel metal2 382398 704 382398 704 0 la_data_out[72]
rlabel metal2 385986 738 385986 738 0 la_data_out[73]
rlabel metal2 389482 840 389482 840 0 la_data_out[74]
rlabel metal2 393070 738 393070 738 0 la_data_out[75]
rlabel metal2 392702 1989 392702 1989 0 la_data_out[76]
rlabel metal2 400154 602 400154 602 0 la_data_out[77]
rlabel metal2 403650 840 403650 840 0 la_data_out[78]
rlabel metal2 407238 806 407238 806 0 la_data_out[79]
rlabel metal2 151846 2047 151846 2047 0 la_data_out[7]
rlabel metal2 410826 602 410826 602 0 la_data_out[80]
rlabel metal2 410090 2499 410090 2499 0 la_data_out[81]
rlabel metal2 417910 772 417910 772 0 la_data_out[82]
rlabel metal2 421406 602 421406 602 0 la_data_out[83]
rlabel metal2 424994 738 424994 738 0 la_data_out[84]
rlabel metal2 428490 806 428490 806 0 la_data_out[85]
rlabel metal2 431894 833 431894 833 0 la_data_out[86]
rlabel metal2 431066 1921 431066 1921 0 la_data_out[87]
rlabel metal2 439162 568 439162 568 0 la_data_out[88]
rlabel metal2 442658 636 442658 636 0 la_data_out[89]
rlabel metal2 155671 340 155671 340 0 la_data_out[8]
rlabel metal2 446055 340 446055 340 0 la_data_out[90]
rlabel metal2 449834 806 449834 806 0 la_data_out[91]
rlabel metal2 448454 2533 448454 2533 0 la_data_out[92]
rlabel metal2 456727 340 456727 340 0 la_data_out[93]
rlabel metal2 460269 340 460269 340 0 la_data_out[94]
rlabel metal2 464002 840 464002 840 0 la_data_out[95]
rlabel metal2 467498 806 467498 806 0 la_data_out[96]
rlabel metal2 465842 2465 465842 2465 0 la_data_out[97]
rlabel metal2 469338 1989 469338 1989 0 la_data_out[98]
rlabel metal2 478170 738 478170 738 0 la_data_out[99]
rlabel metal2 159167 340 159167 340 0 la_data_out[9]
rlabel metal2 128202 806 128202 806 0 la_oenb[0]
rlabel metal2 482671 340 482671 340 0 la_oenb[100]
rlabel metal2 486450 840 486450 840 0 la_oenb[101]
rlabel metal2 484334 2363 484334 2363 0 la_oenb[102]
rlabel metal2 487830 2533 487830 2533 0 la_oenb[103]
rlabel metal2 497122 636 497122 636 0 la_oenb[104]
rlabel metal2 500618 704 500618 704 0 la_oenb[105]
rlabel metal2 504015 340 504015 340 0 la_oenb[106]
rlabel metal2 507511 340 507511 340 0 la_oenb[107]
rlabel metal2 505218 2465 505218 2465 0 la_oenb[108]
rlabel metal2 508714 1989 508714 1989 0 la_oenb[109]
rlabel metal2 163905 340 163905 340 0 la_oenb[10]
rlabel metal2 518183 340 518183 340 0 la_oenb[110]
rlabel via1 521686 85 521686 85 0 la_oenb[111]
rlabel metal2 525458 840 525458 840 0 la_oenb[112]
rlabel metal2 522698 2465 522698 2465 0 la_oenb[113]
rlabel metal2 526102 2533 526102 2533 0 la_oenb[114]
rlabel metal2 536130 704 536130 704 0 la_oenb[115]
rlabel metal2 539626 670 539626 670 0 la_oenb[116]
rlabel metal2 543023 340 543023 340 0 la_oenb[117]
rlabel metal2 546710 772 546710 772 0 la_oenb[118]
rlabel metal2 543490 2499 543490 2499 0 la_oenb[119]
rlabel metal2 167401 340 167401 340 0 la_oenb[11]
rlabel metal2 546986 2057 546986 2057 0 la_oenb[120]
rlabel metal2 557382 806 557382 806 0 la_oenb[121]
rlabel metal2 560878 466 560878 466 0 la_oenb[122]
rlabel metal2 564466 534 564466 534 0 la_oenb[123]
rlabel metal2 560970 2533 560970 2533 0 la_oenb[124]
rlabel metal2 564282 1955 564282 1955 0 la_oenb[125]
rlabel metal2 575138 738 575138 738 0 la_oenb[126]
rlabel metal2 578634 840 578634 840 0 la_oenb[127]
rlabel metal2 170798 2047 170798 2047 0 la_oenb[12]
rlabel metal2 174294 2047 174294 2047 0 la_oenb[13]
rlabel metal2 177981 340 177981 340 0 la_oenb[14]
rlabel metal2 181470 2047 181470 2047 0 la_oenb[15]
rlabel metal2 184966 2047 184966 2047 0 la_oenb[16]
rlabel metal2 188554 2047 188554 2047 0 la_oenb[17]
rlabel metal2 192050 2047 192050 2047 0 la_oenb[18]
rlabel metal2 195539 204 195539 204 0 la_oenb[19]
rlabel metal2 132802 2533 132802 2533 0 la_oenb[1]
rlabel metal2 199035 204 199035 204 0 la_oenb[20]
rlabel metal2 202722 2047 202722 2047 0 la_oenb[21]
rlabel metal2 206218 2047 206218 2047 0 la_oenb[22]
rlabel metal2 209776 340 209776 340 0 la_oenb[23]
rlabel metal2 213394 2047 213394 2047 0 la_oenb[24]
rlabel metal2 216890 2064 216890 2064 0 la_oenb[25]
rlabel metal2 220241 340 220241 340 0 la_oenb[26]
rlabel metal2 223737 340 223737 340 0 la_oenb[27]
rlabel metal2 227562 2047 227562 2047 0 la_oenb[28]
rlabel metal2 231058 2064 231058 2064 0 la_oenb[29]
rlabel metal2 135286 2047 135286 2047 0 la_oenb[2]
rlabel metal2 234646 2064 234646 2064 0 la_oenb[30]
rlabel metal2 238142 2064 238142 2064 0 la_oenb[31]
rlabel metal2 241730 2064 241730 2064 0 la_oenb[32]
rlabel metal2 245226 2098 245226 2098 0 la_oenb[33]
rlabel metal2 248715 340 248715 340 0 la_oenb[34]
rlabel metal2 252402 1588 252402 1588 0 la_oenb[35]
rlabel metal2 255898 1588 255898 1588 0 la_oenb[36]
rlabel metal2 259486 2064 259486 2064 0 la_oenb[37]
rlabel metal2 262982 2098 262982 2098 0 la_oenb[38]
rlabel metal2 266570 2064 266570 2064 0 la_oenb[39]
rlabel metal2 138874 806 138874 806 0 la_oenb[3]
rlabel metal2 270066 2098 270066 2098 0 la_oenb[40]
rlabel metal2 273654 2064 273654 2064 0 la_oenb[41]
rlabel metal2 277150 2098 277150 2098 0 la_oenb[42]
rlabel metal2 280738 2064 280738 2064 0 la_oenb[43]
rlabel metal2 284326 840 284326 840 0 la_oenb[44]
rlabel metal2 287822 2132 287822 2132 0 la_oenb[45]
rlabel metal2 291410 806 291410 806 0 la_oenb[46]
rlabel metal2 294906 2098 294906 2098 0 la_oenb[47]
rlabel metal2 296470 2499 296470 2499 0 la_oenb[48]
rlabel metal2 301990 2098 301990 2098 0 la_oenb[49]
rlabel metal2 142462 2047 142462 2047 0 la_oenb[4]
rlabel metal2 305578 806 305578 806 0 la_oenb[50]
rlabel metal2 309074 2098 309074 2098 0 la_oenb[51]
rlabel metal2 312662 840 312662 840 0 la_oenb[52]
rlabel metal2 313858 2533 313858 2533 0 la_oenb[53]
rlabel metal2 319746 840 319746 840 0 la_oenb[54]
rlabel metal2 323334 738 323334 738 0 la_oenb[55]
rlabel metal2 326830 806 326830 806 0 la_oenb[56]
rlabel metal2 330418 738 330418 738 0 la_oenb[57]
rlabel metal2 333914 772 333914 772 0 la_oenb[58]
rlabel metal2 334742 2499 334742 2499 0 la_oenb[59]
rlabel metal2 145958 840 145958 840 0 la_oenb[5]
rlabel metal2 340998 534 340998 534 0 la_oenb[60]
rlabel metal2 344586 772 344586 772 0 la_oenb[61]
rlabel metal2 348082 840 348082 840 0 la_oenb[62]
rlabel metal2 351670 806 351670 806 0 la_oenb[63]
rlabel metal2 352130 2499 352130 2499 0 la_oenb[64]
rlabel metal2 358754 806 358754 806 0 la_oenb[65]
rlabel metal2 362342 806 362342 806 0 la_oenb[66]
rlabel metal2 365838 840 365838 840 0 la_oenb[67]
rlabel metal2 369426 534 369426 534 0 la_oenb[68]
rlabel metal2 372922 534 372922 534 0 la_oenb[69]
rlabel metal2 149783 340 149783 340 0 la_oenb[6]
rlabel metal2 373014 2499 373014 2499 0 la_oenb[70]
rlabel metal2 380006 840 380006 840 0 la_oenb[71]
rlabel metal2 383594 670 383594 670 0 la_oenb[72]
rlabel metal2 386991 340 386991 340 0 la_oenb[73]
rlabel metal2 390678 704 390678 704 0 la_oenb[74]
rlabel metal2 390402 2465 390402 2465 0 la_oenb[75]
rlabel metal2 397762 806 397762 806 0 la_oenb[76]
rlabel metal2 401350 738 401350 738 0 la_oenb[77]
rlabel metal2 404846 772 404846 772 0 la_oenb[78]
rlabel metal2 408434 738 408434 738 0 la_oenb[79]
rlabel metal2 153279 340 153279 340 0 la_oenb[7]
rlabel metal2 411930 772 411930 772 0 la_oenb[80]
rlabel metal2 411194 3281 411194 3281 0 la_oenb[81]
rlabel metal2 419014 670 419014 670 0 la_oenb[82]
rlabel metal2 422602 806 422602 806 0 la_oenb[83]
rlabel via1 425822 221 425822 221 0 la_oenb[84]
rlabel metal2 429686 704 429686 704 0 la_oenb[85]
rlabel metal2 428674 2431 428674 2431 0 la_oenb[86]
rlabel metal2 436770 670 436770 670 0 la_oenb[87]
rlabel metal2 440167 340 440167 340 0 la_oenb[88]
rlabel metal2 443854 704 443854 704 0 la_oenb[89]
rlabel metal2 156630 2047 156630 2047 0 la_oenb[8]
rlabel metal2 447442 840 447442 840 0 la_oenb[90]
rlabel metal2 450938 772 450938 772 0 la_oenb[91]
rlabel metal2 449558 3281 449558 3281 0 la_oenb[92]
rlabel metal2 458114 670 458114 670 0 la_oenb[93]
rlabel metal2 461610 806 461610 806 0 la_oenb[94]
rlabel via1 465014 85 465014 85 0 la_oenb[95]
rlabel metal2 468694 602 468694 602 0 la_oenb[96]
rlabel metal2 466946 2397 466946 2397 0 la_oenb[97]
rlabel metal2 470442 1921 470442 1921 0 la_oenb[98]
rlabel metal2 479366 670 479366 670 0 la_oenb[99]
rlabel metal2 160126 2047 160126 2047 0 la_oenb[9]
rlabel via1 579646 51 579646 51 0 user_clock2
rlabel via1 581210 323 581210 323 0 user_irq[0]
rlabel via1 581854 187 581854 187 0 user_irq[1]
rlabel via1 583602 85 583602 85 0 user_irq[2]
rlabel metal2 598 2064 598 2064 0 wb_clk_i
rlabel metal2 1702 2098 1702 2098 0 wb_rst_i
rlabel metal2 3089 340 3089 340 0 wbs_ack_o
rlabel metal2 7682 2064 7682 2064 0 wbs_adr_i[0]
rlabel metal2 47886 2064 47886 2064 0 wbs_adr_i[10]
rlabel metal2 51382 2064 51382 2064 0 wbs_adr_i[11]
rlabel metal2 57406 3886 57406 3886 0 wbs_adr_i[12]
rlabel metal2 58466 2064 58466 2064 0 wbs_adr_i[13]
rlabel metal2 62054 1588 62054 1588 0 wbs_adr_i[14]
rlabel metal2 65550 1588 65550 1588 0 wbs_adr_i[15]
rlabel metal2 69138 466 69138 466 0 wbs_adr_i[16]
rlabel metal2 74886 3954 74886 3954 0 wbs_adr_i[17]
rlabel metal2 76222 840 76222 840 0 wbs_adr_i[18]
rlabel metal2 79718 2064 79718 2064 0 wbs_adr_i[19]
rlabel metal2 12374 2064 12374 2064 0 wbs_adr_i[1]
rlabel metal2 83306 840 83306 840 0 wbs_adr_i[20]
rlabel metal2 86894 2064 86894 2064 0 wbs_adr_i[21]
rlabel metal2 90390 806 90390 806 0 wbs_adr_i[22]
rlabel metal2 93978 840 93978 840 0 wbs_adr_i[23]
rlabel metal2 97474 840 97474 840 0 wbs_adr_i[24]
rlabel metal2 101062 840 101062 840 0 wbs_adr_i[25]
rlabel metal2 104558 840 104558 840 0 wbs_adr_i[26]
rlabel metal2 108146 806 108146 806 0 wbs_adr_i[27]
rlabel metal2 111642 738 111642 738 0 wbs_adr_i[28]
rlabel metal2 115230 806 115230 806 0 wbs_adr_i[29]
rlabel metal2 17066 1588 17066 1588 0 wbs_adr_i[2]
rlabel metal2 119055 340 119055 340 0 wbs_adr_i[30]
rlabel metal2 122314 806 122314 806 0 wbs_adr_i[31]
rlabel metal2 21850 2064 21850 2064 0 wbs_adr_i[3]
rlabel metal2 26542 2098 26542 2098 0 wbs_adr_i[4]
rlabel metal2 30130 2098 30130 2098 0 wbs_adr_i[5]
rlabel metal2 36614 3920 36614 3920 0 wbs_adr_i[6]
rlabel metal2 37214 2098 37214 2098 0 wbs_adr_i[7]
rlabel metal2 40710 2064 40710 2064 0 wbs_adr_i[8]
rlabel metal2 44298 2064 44298 2064 0 wbs_adr_i[9]
rlabel metal2 4094 1588 4094 1588 0 wbs_cyc_i
rlabel metal2 8786 636 8786 636 0 wbs_dat_i[0]
rlabel metal2 48990 2098 48990 2098 0 wbs_dat_i[10]
rlabel metal2 52578 534 52578 534 0 wbs_dat_i[11]
rlabel metal2 56074 2132 56074 2132 0 wbs_dat_i[12]
rlabel metal2 59662 534 59662 534 0 wbs_dat_i[13]
rlabel metal2 63250 1690 63250 1690 0 wbs_dat_i[14]
rlabel metal2 66937 340 66937 340 0 wbs_dat_i[15]
rlabel metal2 70334 2064 70334 2064 0 wbs_dat_i[16]
rlabel metal2 75990 3886 75990 3886 0 wbs_dat_i[17]
rlabel metal2 77418 806 77418 806 0 wbs_dat_i[18]
rlabel metal2 80914 2098 80914 2098 0 wbs_dat_i[19]
rlabel metal2 16834 3920 16834 3920 0 wbs_dat_i[1]
rlabel metal2 84502 806 84502 806 0 wbs_dat_i[20]
rlabel metal2 87998 2098 87998 2098 0 wbs_dat_i[21]
rlabel metal2 91586 840 91586 840 0 wbs_dat_i[22]
rlabel metal2 95174 2064 95174 2064 0 wbs_dat_i[23]
rlabel metal2 98670 806 98670 806 0 wbs_dat_i[24]
rlabel metal2 102258 806 102258 806 0 wbs_dat_i[25]
rlabel metal2 105754 534 105754 534 0 wbs_dat_i[26]
rlabel metal2 109342 840 109342 840 0 wbs_dat_i[27]
rlabel metal2 114218 2533 114218 2533 0 wbs_dat_i[28]
rlabel metal2 116426 840 116426 840 0 wbs_dat_i[29]
rlabel metal2 18262 1622 18262 1622 0 wbs_dat_i[2]
rlabel metal2 119922 840 119922 840 0 wbs_dat_i[30]
rlabel metal2 123510 738 123510 738 0 wbs_dat_i[31]
rlabel metal2 23046 2098 23046 2098 0 wbs_dat_i[3]
rlabel metal2 27738 2132 27738 2132 0 wbs_dat_i[4]
rlabel metal2 31326 2064 31326 2064 0 wbs_dat_i[5]
rlabel metal2 37718 3886 37718 3886 0 wbs_dat_i[6]
rlabel metal2 38410 2132 38410 2132 0 wbs_dat_i[7]
rlabel metal2 41906 2098 41906 2098 0 wbs_dat_i[8]
rlabel metal2 45494 2098 45494 2098 0 wbs_dat_i[9]
rlabel metal2 9982 1588 9982 1588 0 wbs_dat_o[0]
rlabel metal2 50186 2132 50186 2132 0 wbs_dat_o[10]
rlabel metal2 56302 3920 56302 3920 0 wbs_dat_o[11]
rlabel metal2 57270 2098 57270 2098 0 wbs_dat_o[12]
rlabel metal2 60858 840 60858 840 0 wbs_dat_o[13]
rlabel metal2 64354 2064 64354 2064 0 wbs_dat_o[14]
rlabel metal2 67942 840 67942 840 0 wbs_dat_o[15]
rlabel metal2 71530 2098 71530 2098 0 wbs_dat_o[16]
rlabel metal2 75026 806 75026 806 0 wbs_dat_o[17]
rlabel metal2 78614 2098 78614 2098 0 wbs_dat_o[18]
rlabel metal2 82110 806 82110 806 0 wbs_dat_o[19]
rlabel metal2 18030 3954 18030 3954 0 wbs_dat_o[1]
rlabel metal2 85698 840 85698 840 0 wbs_dat_o[20]
rlabel metal2 89194 840 89194 840 0 wbs_dat_o[21]
rlabel metal2 94530 2499 94530 2499 0 wbs_dat_o[22]
rlabel metal2 96278 2098 96278 2098 0 wbs_dat_o[23]
rlabel metal2 99866 772 99866 772 0 wbs_dat_o[24]
rlabel metal2 103362 2064 103362 2064 0 wbs_dat_o[25]
rlabel metal2 106950 840 106950 840 0 wbs_dat_o[26]
rlabel metal2 110538 806 110538 806 0 wbs_dat_o[27]
rlabel metal2 114034 772 114034 772 0 wbs_dat_o[28]
rlabel metal2 117622 806 117622 806 0 wbs_dat_o[29]
rlabel metal2 19458 2098 19458 2098 0 wbs_dat_o[2]
rlabel metal2 121118 636 121118 636 0 wbs_dat_o[30]
rlabel metal2 124706 806 124706 806 0 wbs_dat_o[31]
rlabel metal2 24242 2132 24242 2132 0 wbs_dat_o[3]
rlabel metal2 28934 1588 28934 1588 0 wbs_dat_o[4]
rlabel metal2 32430 2132 32430 2132 0 wbs_dat_o[5]
rlabel metal2 36018 1588 36018 1588 0 wbs_dat_o[6]
rlabel metal2 39606 1588 39606 1588 0 wbs_dat_o[7]
rlabel metal2 43102 2132 43102 2132 0 wbs_dat_o[8]
rlabel metal2 46690 2132 46690 2132 0 wbs_dat_o[9]
rlabel metal2 11178 2132 11178 2132 0 wbs_sel_i[0]
rlabel metal2 19134 3886 19134 3886 0 wbs_sel_i[1]
rlabel metal2 20654 2132 20654 2132 0 wbs_sel_i[2]
rlabel metal2 25346 2064 25346 2064 0 wbs_sel_i[3]
rlabel metal2 5481 340 5481 340 0 wbs_stb_i
rlabel metal2 6486 1690 6486 1690 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
